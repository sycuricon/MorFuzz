module IntXbar(
  input         auto_int_in_0,
  output        auto_int_out_0,
  output [29:0] io_covSum
);
  wire [29:0] IntXbar_covSum;
  assign auto_int_out_0 = auto_int_in_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign IntXbar_covSum = 30'h0;
  assign io_covSum = IntXbar_covSum;
endmodule
module SimpleClockGroupSource(
  input         clock,
  input         reset,
  output        auto_out_member_subsystem_sbus_5_clock,
  output        auto_out_member_subsystem_sbus_5_reset,
  output        auto_out_member_subsystem_sbus_4_clock,
  output        auto_out_member_subsystem_sbus_4_reset,
  output        auto_out_member_subsystem_sbus_3_clock,
  output        auto_out_member_subsystem_sbus_3_reset,
  output        auto_out_member_subsystem_sbus_2_clock,
  output        auto_out_member_subsystem_sbus_2_reset,
  output        auto_out_member_subsystem_sbus_1_clock,
  output        auto_out_member_subsystem_sbus_1_reset,
  output        auto_out_member_subsystem_sbus_0_clock,
  output        auto_out_member_subsystem_sbus_0_reset,
  output [29:0] io_covSum
);
  wire [29:0] SimpleClockGroupSource_covSum;
  assign auto_out_member_subsystem_sbus_5_clock = clock; // @[Nodes.scala 1207:84 ClockGroup.scala 72:17]
  assign auto_out_member_subsystem_sbus_5_reset = reset; // @[Nodes.scala 1207:84 ClockGroup.scala 72:35]
  assign auto_out_member_subsystem_sbus_4_clock = clock; // @[Nodes.scala 1207:84 ClockGroup.scala 72:17]
  assign auto_out_member_subsystem_sbus_4_reset = reset; // @[Nodes.scala 1207:84 ClockGroup.scala 72:35]
  assign auto_out_member_subsystem_sbus_3_clock = clock; // @[Nodes.scala 1207:84 ClockGroup.scala 72:17]
  assign auto_out_member_subsystem_sbus_3_reset = reset; // @[Nodes.scala 1207:84 ClockGroup.scala 72:35]
  assign auto_out_member_subsystem_sbus_2_clock = clock; // @[Nodes.scala 1207:84 ClockGroup.scala 72:17]
  assign auto_out_member_subsystem_sbus_2_reset = reset; // @[Nodes.scala 1207:84 ClockGroup.scala 72:35]
  assign auto_out_member_subsystem_sbus_1_clock = clock; // @[Nodes.scala 1207:84 ClockGroup.scala 72:17]
  assign auto_out_member_subsystem_sbus_1_reset = reset; // @[Nodes.scala 1207:84 ClockGroup.scala 72:35]
  assign auto_out_member_subsystem_sbus_0_clock = clock; // @[Nodes.scala 1207:84 ClockGroup.scala 72:17]
  assign auto_out_member_subsystem_sbus_0_reset = reset; // @[Nodes.scala 1207:84 ClockGroup.scala 72:35]
  assign SimpleClockGroupSource_covSum = 30'h0;
  assign io_covSum = SimpleClockGroupSource_covSum;
endmodule
module FixedClockBroadcast(
  input         auto_in_clock,
  input         auto_in_reset,
  output        auto_out_2_clock,
  output        auto_out_2_reset,
  output        auto_out_1_clock,
  output        auto_out_1_reset,
  output        auto_out_0_clock,
  output        auto_out_0_reset,
  output [29:0] io_covSum
);
  wire [29:0] FixedClockBroadcast_covSum;
  assign auto_out_2_clock = auto_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_2_reset = auto_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_clock = auto_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_reset = auto_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_clock = auto_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_reset = auto_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign FixedClockBroadcast_covSum = 30'h0;
  assign io_covSum = FixedClockBroadcast_covSum;
endmodule
module TLXbar(
  input         clock,
  input         reset,
  output        auto_in_1_a_ready,
  input         auto_in_1_a_valid,
  input  [2:0]  auto_in_1_a_bits_opcode,
  input  [2:0]  auto_in_1_a_bits_param,
  input  [3:0]  auto_in_1_a_bits_size,
  input  [5:0]  auto_in_1_a_bits_source,
  input  [31:0] auto_in_1_a_bits_address,
  input         auto_in_1_a_bits_user_amba_prot_bufferable,
  input         auto_in_1_a_bits_user_amba_prot_modifiable,
  input         auto_in_1_a_bits_user_amba_prot_readalloc,
  input         auto_in_1_a_bits_user_amba_prot_writealloc,
  input         auto_in_1_a_bits_user_amba_prot_privileged,
  input         auto_in_1_a_bits_user_amba_prot_secure,
  input         auto_in_1_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_1_a_bits_mask,
  input  [63:0] auto_in_1_a_bits_data,
  input         auto_in_1_d_ready,
  output        auto_in_1_d_valid,
  output [2:0]  auto_in_1_d_bits_opcode,
  output [3:0]  auto_in_1_d_bits_size,
  output [5:0]  auto_in_1_d_bits_source,
  output        auto_in_1_d_bits_denied,
  output [63:0] auto_in_1_d_bits_data,
  output        auto_in_1_d_bits_corrupt,
  output        auto_in_0_a_ready,
  input         auto_in_0_a_valid,
  input  [2:0]  auto_in_0_a_bits_opcode,
  input  [2:0]  auto_in_0_a_bits_param,
  input  [3:0]  auto_in_0_a_bits_size,
  input  [3:0]  auto_in_0_a_bits_source,
  input  [31:0] auto_in_0_a_bits_address,
  input         auto_in_0_a_bits_user_amba_prot_bufferable,
  input         auto_in_0_a_bits_user_amba_prot_modifiable,
  input         auto_in_0_a_bits_user_amba_prot_readalloc,
  input         auto_in_0_a_bits_user_amba_prot_writealloc,
  input         auto_in_0_a_bits_user_amba_prot_privileged,
  input         auto_in_0_a_bits_user_amba_prot_secure,
  input         auto_in_0_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_0_a_bits_mask,
  input  [63:0] auto_in_0_a_bits_data,
  input         auto_in_0_d_ready,
  output        auto_in_0_d_valid,
  output [2:0]  auto_in_0_d_bits_opcode,
  output [3:0]  auto_in_0_d_bits_size,
  output [3:0]  auto_in_0_d_bits_source,
  output        auto_in_0_d_bits_denied,
  output [63:0] auto_in_0_d_bits_data,
  output        auto_in_0_d_bits_corrupt,
  input         auto_out_1_a_ready,
  output        auto_out_1_a_valid,
  output [2:0]  auto_out_1_a_bits_opcode,
  output [2:0]  auto_out_1_a_bits_size,
  output [6:0]  auto_out_1_a_bits_source,
  output [31:0] auto_out_1_a_bits_address,
  output        auto_out_1_a_bits_user_amba_prot_bufferable,
  output        auto_out_1_a_bits_user_amba_prot_modifiable,
  output        auto_out_1_a_bits_user_amba_prot_readalloc,
  output        auto_out_1_a_bits_user_amba_prot_writealloc,
  output        auto_out_1_a_bits_user_amba_prot_privileged,
  output        auto_out_1_a_bits_user_amba_prot_secure,
  output        auto_out_1_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_1_a_bits_mask,
  output [63:0] auto_out_1_a_bits_data,
  output        auto_out_1_d_ready,
  input         auto_out_1_d_valid,
  input  [2:0]  auto_out_1_d_bits_opcode,
  input  [2:0]  auto_out_1_d_bits_size,
  input  [6:0]  auto_out_1_d_bits_source,
  input         auto_out_1_d_bits_denied,
  input  [63:0] auto_out_1_d_bits_data,
  input         auto_out_1_d_bits_corrupt,
  input         auto_out_0_a_ready,
  output        auto_out_0_a_valid,
  output [2:0]  auto_out_0_a_bits_opcode,
  output [2:0]  auto_out_0_a_bits_param,
  output [3:0]  auto_out_0_a_bits_size,
  output [6:0]  auto_out_0_a_bits_source,
  output [30:0] auto_out_0_a_bits_address,
  output [7:0]  auto_out_0_a_bits_mask,
  output [63:0] auto_out_0_a_bits_data,
  output        auto_out_0_d_ready,
  input         auto_out_0_d_valid,
  input  [2:0]  auto_out_0_d_bits_opcode,
  input  [3:0]  auto_out_0_d_bits_size,
  input  [6:0]  auto_out_0_d_bits_source,
  input         auto_out_0_d_bits_denied,
  input  [63:0] auto_out_0_d_bits_data,
  input         auto_out_0_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] _GEN_4 = {{3'd0}, auto_in_0_a_bits_source}; // @[Xbar.scala 237:55]
  wire [6:0] in_0_a_bits_source = _GEN_4 | 7'h40; // @[Xbar.scala 237:55]
  reg [8:0] beatsLeft_2; // @[Arbiter.scala 87:30]
  wire  idle_2 = beatsLeft_2 == 9'h0; // @[Arbiter.scala 88:28]
  wire  requestDOI_1_0 = auto_out_1_d_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  portsDIO_filtered_1_0_valid = auto_out_1_d_valid & requestDOI_1_0; // @[Xbar.scala 179:40]
  wire  requestDOI_0_0 = auto_out_0_d_bits_source[6:4] == 3'h4; // @[Parameters.scala 54:32]
  wire  portsDIO_filtered__0_valid = auto_out_0_d_valid & requestDOI_0_0; // @[Xbar.scala 179:40]
  wire [1:0] readys_valid_2 = {portsDIO_filtered_1_0_valid,portsDIO_filtered__0_valid}; // @[Cat.scala 31:58]
  reg [1:0] readys_mask_2; // @[Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T_4 = ~readys_mask_2; // @[Arbiter.scala 24:30]
  wire [1:0] _readys_filter_T_5 = readys_valid_2 & _readys_filter_T_4; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter_2 = {_readys_filter_T_5,portsDIO_filtered_1_0_valid,portsDIO_filtered__0_valid}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_5 = {{1'd0}, readys_filter_2[3:1]}; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_11 = readys_filter_2 | _GEN_5; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_14 = {readys_mask_2, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_6 = {{1'd0}, _readys_unready_T_11[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready_2 = _GEN_6 | _readys_unready_T_14; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_8 = readys_unready_2[3:2] & readys_unready_2[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys_2 = ~_readys_readys_T_8; // @[Arbiter.scala 26:18]
  wire  readys_2_0 = readys_readys_2[0]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_2_0 = readys_2_0 & portsDIO_filtered__0_valid; // @[Arbiter.scala 97:79]
  reg  state_2_0; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_2_0 = idle_2 ? earlyWinner_2_0 : state_2_0; // @[Arbiter.scala 117:30]
  wire [6:0] _T_174 = muxStateEarly_2_0 ? auto_out_0_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire  readys_2_1 = readys_readys_2[1]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_2_1 = readys_2_1 & portsDIO_filtered_1_0_valid; // @[Arbiter.scala 97:79]
  reg  state_2_1; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_2_1 = idle_2 ? earlyWinner_2_1 : state_2_1; // @[Arbiter.scala 117:30]
  wire [6:0] _T_175 = muxStateEarly_2_1 ? auto_out_1_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] sink_ACancel_5_bits_source = _T_174 | _T_175; // @[Mux.scala 27:73]
  reg [8:0] beatsLeft_3; // @[Arbiter.scala 87:30]
  wire  idle_3 = beatsLeft_3 == 9'h0; // @[Arbiter.scala 88:28]
  wire  requestDOI_1_1 = ~auto_out_1_d_bits_source[6]; // @[Parameters.scala 54:32]
  wire  portsDIO_filtered_1_1_valid = auto_out_1_d_valid & requestDOI_1_1; // @[Xbar.scala 179:40]
  wire  requestDOI_0_1 = ~auto_out_0_d_bits_source[6]; // @[Parameters.scala 54:32]
  wire  portsDIO_filtered__1_valid = auto_out_0_d_valid & requestDOI_0_1; // @[Xbar.scala 179:40]
  wire [1:0] readys_valid_3 = {portsDIO_filtered_1_1_valid,portsDIO_filtered__1_valid}; // @[Cat.scala 31:58]
  reg [1:0] readys_mask_3; // @[Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T_6 = ~readys_mask_3; // @[Arbiter.scala 24:30]
  wire [1:0] _readys_filter_T_7 = readys_valid_3 & _readys_filter_T_6; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter_3 = {_readys_filter_T_7,portsDIO_filtered_1_1_valid,portsDIO_filtered__1_valid}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_7 = {{1'd0}, readys_filter_3[3:1]}; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_16 = readys_filter_3 | _GEN_7; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_19 = {readys_mask_3, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_8 = {{1'd0}, _readys_unready_T_16[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready_3 = _GEN_8 | _readys_unready_T_19; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_11 = readys_unready_3[3:2] & readys_unready_3[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys_3 = ~_readys_readys_T_11; // @[Arbiter.scala 26:18]
  wire  readys_3_0 = readys_readys_3[0]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_3_0 = readys_3_0 & portsDIO_filtered__1_valid; // @[Arbiter.scala 97:79]
  reg  state_3_0; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_3_0 = idle_3 ? earlyWinner_3_0 : state_3_0; // @[Arbiter.scala 117:30]
  wire [6:0] _T_222 = muxStateEarly_3_0 ? auto_out_0_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire  readys_3_1 = readys_readys_3[1]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_3_1 = readys_3_1 & portsDIO_filtered_1_1_valid; // @[Arbiter.scala 97:79]
  reg  state_3_1; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_3_1 = idle_3 ? earlyWinner_3_1 : state_3_1; // @[Arbiter.scala 117:30]
  wire [6:0] _T_223 = muxStateEarly_3_1 ? auto_out_1_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] sink_ACancel_7_bits_source = _T_222 | _T_223; // @[Mux.scala 27:73]
  wire [32:0] _requestAIO_T_1 = {1'b0,$signed(auto_in_0_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_3 = $signed(_requestAIO_T_1) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_0 = $signed(_requestAIO_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_5 = auto_in_0_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_6 = {1'b0,$signed(_requestAIO_T_5)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_8 = $signed(_requestAIO_T_6) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_1 = $signed(_requestAIO_T_8) == 33'sh0; // @[Parameters.scala 137:67]
  wire [32:0] _requestAIO_T_11 = {1'b0,$signed(auto_in_1_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_13 = $signed(_requestAIO_T_11) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  requestAIO_1_0 = $signed(_requestAIO_T_13) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_15 = auto_in_1_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_16 = {1'b0,$signed(_requestAIO_T_15)}; // @[Parameters.scala 137:49]
  wire [32:0] _requestAIO_T_18 = $signed(_requestAIO_T_16) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  requestAIO_1_1 = $signed(_requestAIO_T_18) == 33'sh0; // @[Parameters.scala 137:67]
  wire [26:0] _beatsAI_decode_T_1 = 27'hfff << auto_in_0_a_bits_size; // @[package.scala 234:77]
  wire [11:0] _beatsAI_decode_T_3 = ~_beatsAI_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] beatsAI_decode = _beatsAI_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  beatsAI_opdata = ~auto_in_0_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [8:0] beatsAI_0 = beatsAI_opdata ? beatsAI_decode : 9'h0; // @[Edges.scala 220:14]
  wire [26:0] _beatsAI_decode_T_5 = 27'hfff << auto_in_1_a_bits_size; // @[package.scala 234:77]
  wire [11:0] _beatsAI_decode_T_7 = ~_beatsAI_decode_T_5[11:0]; // @[package.scala 234:46]
  wire [8:0] beatsAI_decode_1 = _beatsAI_decode_T_7[11:3]; // @[Edges.scala 219:59]
  wire  beatsAI_opdata_1 = ~auto_in_1_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [8:0] beatsAI_1 = beatsAI_opdata_1 ? beatsAI_decode_1 : 9'h0; // @[Edges.scala 220:14]
  wire [26:0] _beatsDO_decode_T_1 = 27'hfff << auto_out_0_d_bits_size; // @[package.scala 234:77]
  wire [11:0] _beatsDO_decode_T_3 = ~_beatsDO_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] beatsDO_decode = _beatsDO_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata = auto_out_0_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [8:0] beatsDO_0 = beatsDO_opdata ? beatsDO_decode : 9'h0; // @[Edges.scala 220:14]
  wire [3:0] out_2_1_d_bits_size = {{1'd0}, auto_out_1_d_bits_size}; // @[BundleMap.scala 247:19 Xbar.scala 288:19]
  wire [20:0] _beatsDO_decode_T_5 = 21'h3f << out_2_1_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_7 = ~_beatsDO_decode_T_5[5:0]; // @[package.scala 234:46]
  wire [2:0] beatsDO_decode_1 = _beatsDO_decode_T_7[5:3]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata_1 = auto_out_1_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] beatsDO_1 = beatsDO_opdata_1 ? beatsDO_decode_1 : 3'h0; // @[Edges.scala 220:14]
  wire  portsAOI_filtered__0_earlyValid = auto_in_0_a_valid & requestAIO_0_0; // @[Xbar.scala 428:50]
  wire  portsAOI_filtered__1_earlyValid = auto_in_0_a_valid & requestAIO_0_1; // @[Xbar.scala 428:50]
  reg [8:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 9'h0; // @[Arbiter.scala 88:28]
  wire  portsAOI_filtered_1_0_earlyValid = auto_in_1_a_valid & requestAIO_1_0; // @[Xbar.scala 428:50]
  wire [1:0] readys_valid = {portsAOI_filtered_1_0_earlyValid,portsAOI_filtered__0_earlyValid}; // @[Cat.scala 31:58]
  reg [1:0] readys_mask; // @[Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 24:30]
  wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter = {_readys_filter_T_1,portsAOI_filtered_1_0_earlyValid,portsAOI_filtered__0_earlyValid}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_9 = {{1'd0}, readys_filter[3:1]}; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_9; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_10 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready = _GEN_10 | _readys_unready_T_4; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 26:18]
  wire  readys__0 = readys_readys[0]; // @[Arbiter.scala 95:86]
  reg  state__0; // @[Arbiter.scala 116:26]
  wire  allowed__0 = idle ? readys__0 : state__0; // @[Arbiter.scala 121:24]
  wire  portsAOI_filtered__0_ready = auto_out_0_a_ready & allowed__0; // @[Arbiter.scala 123:31]
  reg [8:0] beatsLeft_1; // @[Arbiter.scala 87:30]
  wire  idle_1 = beatsLeft_1 == 9'h0; // @[Arbiter.scala 88:28]
  wire  portsAOI_filtered_1_1_earlyValid = auto_in_1_a_valid & requestAIO_1_1; // @[Xbar.scala 428:50]
  wire [1:0] readys_valid_1 = {portsAOI_filtered_1_1_earlyValid,portsAOI_filtered__1_earlyValid}; // @[Cat.scala 31:58]
  reg [1:0] readys_mask_1; // @[Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T_2 = ~readys_mask_1; // @[Arbiter.scala 24:30]
  wire [1:0] _readys_filter_T_3 = readys_valid_1 & _readys_filter_T_2; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter_1 = {_readys_filter_T_3,portsAOI_filtered_1_1_earlyValid,portsAOI_filtered__1_earlyValid}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_11 = {{1'd0}, readys_filter_1[3:1]}; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_6 = readys_filter_1 | _GEN_11; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_9 = {readys_mask_1, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_12 = {{1'd0}, _readys_unready_T_6[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready_1 = _GEN_12 | _readys_unready_T_9; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_5 = readys_unready_1[3:2] & readys_unready_1[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys_1 = ~_readys_readys_T_5; // @[Arbiter.scala 26:18]
  wire  readys_1_0 = readys_readys_1[0]; // @[Arbiter.scala 95:86]
  reg  state_1_0; // @[Arbiter.scala 116:26]
  wire  allowed_1_0 = idle_1 ? readys_1_0 : state_1_0; // @[Arbiter.scala 121:24]
  wire  portsAOI_filtered__1_ready = auto_out_1_a_ready & allowed_1_0; // @[Arbiter.scala 123:31]
  wire  readys__1 = readys_readys[1]; // @[Arbiter.scala 95:86]
  reg  state__1; // @[Arbiter.scala 116:26]
  wire  allowed__1 = idle ? readys__1 : state__1; // @[Arbiter.scala 121:24]
  wire  portsAOI_filtered_1_0_ready = auto_out_0_a_ready & allowed__1; // @[Arbiter.scala 123:31]
  wire  readys_1_1 = readys_readys_1[1]; // @[Arbiter.scala 95:86]
  reg  state_1_1; // @[Arbiter.scala 116:26]
  wire  allowed_1_1 = idle_1 ? readys_1_1 : state_1_1; // @[Arbiter.scala 121:24]
  wire  portsAOI_filtered_1_1_ready = auto_out_1_a_ready & allowed_1_1; // @[Arbiter.scala 123:31]
  wire  allowed_2_0 = idle_2 ? readys_2_0 : state_2_0; // @[Arbiter.scala 121:24]
  wire  out_8_ready = auto_in_0_d_ready & allowed_2_0; // @[Arbiter.scala 123:31]
  wire  allowed_3_0 = idle_3 ? readys_3_0 : state_3_0; // @[Arbiter.scala 121:24]
  wire  out_12_ready = auto_in_1_d_ready & allowed_3_0; // @[Arbiter.scala 123:31]
  wire  allowed_2_1 = idle_2 ? readys_2_1 : state_2_1; // @[Arbiter.scala 121:24]
  wire  out_9_ready = auto_in_0_d_ready & allowed_2_1; // @[Arbiter.scala 123:31]
  wire  allowed_3_1 = idle_3 ? readys_3_1 : state_3_1; // @[Arbiter.scala 121:24]
  wire  out_13_ready = auto_in_1_d_ready & allowed_3_1; // @[Arbiter.scala 123:31]
  wire  latch = idle & auto_out_0_a_ready; // @[Arbiter.scala 89:24]
  wire  _readys_T_3 = ~reset; // @[Arbiter.scala 22:12]
  wire [1:0] _readys_mask_T = readys_readys & readys_valid; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[package.scala 244:43]
  wire  earlyWinner__0 = readys__0 & portsAOI_filtered__0_earlyValid; // @[Arbiter.scala 97:79]
  wire  earlyWinner__1 = readys__1 & portsAOI_filtered_1_0_earlyValid; // @[Arbiter.scala 97:79]
  wire  _T_10 = portsAOI_filtered__0_earlyValid | portsAOI_filtered_1_0_earlyValid; // @[Arbiter.scala 107:36]
  wire  _T_11 = ~(portsAOI_filtered__0_earlyValid | portsAOI_filtered_1_0_earlyValid); // @[Arbiter.scala 107:15]
  wire [8:0] maskedBeats_0 = earlyWinner__0 ? beatsAI_0 : 9'h0; // @[Arbiter.scala 111:73]
  wire [8:0] maskedBeats_1 = earlyWinner__1 ? beatsAI_1 : 9'h0; // @[Arbiter.scala 111:73]
  wire [8:0] initBeats = maskedBeats_0 | maskedBeats_1; // @[Arbiter.scala 112:44]
  wire  muxStateEarly__0 = idle ? earlyWinner__0 : state__0; // @[Arbiter.scala 117:30]
  wire  muxStateEarly__1 = idle ? earlyWinner__1 : state__1; // @[Arbiter.scala 117:30]
  wire  _out_0_a_earlyValid_T_3 = state__0 & portsAOI_filtered__0_earlyValid | state__1 &
    portsAOI_filtered_1_0_earlyValid; // @[Mux.scala 27:73]
  wire  out_2_0_a_earlyValid = idle ? _T_10 : _out_0_a_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_out_0_a_ready & out_2_0_a_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [8:0] _GEN_13 = {{8'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [8:0] _beatsLeft_T_4 = beatsLeft - _GEN_13; // @[Arbiter.scala 113:52]
  wire [63:0] _T_27 = muxStateEarly__0 ? auto_in_0_a_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_28 = muxStateEarly__1 ? auto_in_1_a_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_30 = muxStateEarly__0 ? auto_in_0_a_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_31 = muxStateEarly__1 ? auto_in_1_a_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_54 = muxStateEarly__0 ? auto_in_0_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_55 = muxStateEarly__1 ? auto_in_1_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] out_2_0_a_bits_address = _T_54 | _T_55; // @[Mux.scala 27:73]
  wire [6:0] _T_57 = muxStateEarly__0 ? in_0_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] in_1_a_bits_source = {{1'd0}, auto_in_1_a_bits_source}; // @[Xbar.scala 231:18 237:29]
  wire [6:0] _T_58 = muxStateEarly__1 ? in_1_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_60 = muxStateEarly__0 ? auto_in_0_a_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_61 = muxStateEarly__1 ? auto_in_1_a_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_63 = muxStateEarly__0 ? auto_in_0_a_bits_param : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_64 = muxStateEarly__1 ? auto_in_1_a_bits_param : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_66 = muxStateEarly__0 ? auto_in_0_a_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_67 = muxStateEarly__1 ? auto_in_1_a_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire  latch_1 = idle_1 & auto_out_1_a_ready; // @[Arbiter.scala 89:24]
  wire [1:0] _readys_mask_T_5 = readys_readys_1 & readys_valid_1; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_6 = {_readys_mask_T_5, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_8 = _readys_mask_T_5 | _readys_mask_T_6[1:0]; // @[package.scala 244:43]
  wire  earlyWinner_1_0 = readys_1_0 & portsAOI_filtered__1_earlyValid; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1_1 = readys_1_1 & portsAOI_filtered_1_1_earlyValid; // @[Arbiter.scala 97:79]
  wire  _T_79 = portsAOI_filtered__1_earlyValid | portsAOI_filtered_1_1_earlyValid; // @[Arbiter.scala 107:36]
  wire  _T_80 = ~(portsAOI_filtered__1_earlyValid | portsAOI_filtered_1_1_earlyValid); // @[Arbiter.scala 107:15]
  wire [8:0] maskedBeats_0_1 = earlyWinner_1_0 ? beatsAI_0 : 9'h0; // @[Arbiter.scala 111:73]
  wire [8:0] maskedBeats_1_1 = earlyWinner_1_1 ? beatsAI_1 : 9'h0; // @[Arbiter.scala 111:73]
  wire [8:0] initBeats_1 = maskedBeats_0_1 | maskedBeats_1_1; // @[Arbiter.scala 112:44]
  wire  muxStateEarly_1_0 = idle_1 ? earlyWinner_1_0 : state_1_0; // @[Arbiter.scala 117:30]
  wire  muxStateEarly_1_1 = idle_1 ? earlyWinner_1_1 : state_1_1; // @[Arbiter.scala 117:30]
  wire  _out_1_a_earlyValid_T_3 = state_1_0 & portsAOI_filtered__1_earlyValid | state_1_1 &
    portsAOI_filtered_1_1_earlyValid; // @[Mux.scala 27:73]
  wire  out_2_1_a_earlyValid = idle_1 ? _T_79 : _out_1_a_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_8 = auto_out_1_a_ready & out_2_1_a_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [8:0] _GEN_14 = {{8'd0}, _beatsLeft_T_8}; // @[Arbiter.scala 113:52]
  wire [8:0] _beatsLeft_T_10 = beatsLeft_1 - _GEN_14; // @[Arbiter.scala 113:52]
  wire [63:0] _T_96 = muxStateEarly_1_0 ? auto_in_0_a_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_97 = muxStateEarly_1_1 ? auto_in_1_a_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_99 = muxStateEarly_1_0 ? auto_in_0_a_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_100 = muxStateEarly_1_1 ? auto_in_1_a_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_123 = muxStateEarly_1_0 ? auto_in_0_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_124 = muxStateEarly_1_1 ? auto_in_1_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_126 = muxStateEarly_1_0 ? in_0_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_127 = muxStateEarly_1_1 ? in_1_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_129 = muxStateEarly_1_0 ? auto_in_0_a_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_130 = muxStateEarly_1_1 ? auto_in_1_a_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] out_2_1_a_bits_size = _T_129 | _T_130; // @[Mux.scala 27:73]
  wire [2:0] _T_135 = muxStateEarly_1_0 ? auto_in_0_a_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_136 = muxStateEarly_1_1 ? auto_in_1_a_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire  latch_2 = idle_2 & auto_in_0_d_ready; // @[Arbiter.scala 89:24]
  wire [1:0] _readys_mask_T_10 = readys_readys_2 & readys_valid_2; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_11 = {_readys_mask_T_10, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_13 = _readys_mask_T_10 | _readys_mask_T_11[1:0]; // @[package.scala 244:43]
  wire  _T_148 = portsDIO_filtered__0_valid | portsDIO_filtered_1_0_valid; // @[Arbiter.scala 107:36]
  wire  _T_149 = ~(portsDIO_filtered__0_valid | portsDIO_filtered_1_0_valid); // @[Arbiter.scala 107:15]
  wire [8:0] maskedBeats_0_2 = earlyWinner_2_0 ? beatsDO_0 : 9'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_1_2 = earlyWinner_2_1 ? beatsDO_1 : 3'h0; // @[Arbiter.scala 111:73]
  wire [8:0] _GEN_15 = {{6'd0}, maskedBeats_1_2}; // @[Arbiter.scala 112:44]
  wire [8:0] initBeats_2 = maskedBeats_0_2 | _GEN_15; // @[Arbiter.scala 112:44]
  wire  _sink_ACancel_earlyValid_T_3 = state_2_0 & portsDIO_filtered__0_valid | state_2_1 & portsDIO_filtered_1_0_valid; // @[Mux.scala 27:73]
  wire  sink_ACancel_5_earlyValid = idle_2 ? _T_148 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_14 = auto_in_0_d_ready & sink_ACancel_5_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [8:0] _GEN_16 = {{8'd0}, _beatsLeft_T_14}; // @[Arbiter.scala 113:52]
  wire [8:0] _beatsLeft_T_16 = beatsLeft_2 - _GEN_16; // @[Arbiter.scala 113:52]
  wire [63:0] _T_165 = muxStateEarly_2_0 ? auto_out_0_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_166 = muxStateEarly_2_1 ? auto_out_1_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_177 = muxStateEarly_2_0 ? auto_out_0_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_178 = muxStateEarly_2_1 ? out_2_1_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_183 = muxStateEarly_2_0 ? auto_out_0_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_184 = muxStateEarly_2_1 ? auto_out_1_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire  latch_3 = idle_3 & auto_in_1_d_ready; // @[Arbiter.scala 89:24]
  wire [1:0] _readys_mask_T_15 = readys_readys_3 & readys_valid_3; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_16 = {_readys_mask_T_15, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_18 = _readys_mask_T_15 | _readys_mask_T_16[1:0]; // @[package.scala 244:43]
  wire  _T_196 = portsDIO_filtered__1_valid | portsDIO_filtered_1_1_valid; // @[Arbiter.scala 107:36]
  wire  _T_197 = ~(portsDIO_filtered__1_valid | portsDIO_filtered_1_1_valid); // @[Arbiter.scala 107:15]
  wire [8:0] maskedBeats_0_3 = earlyWinner_3_0 ? beatsDO_0 : 9'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_1_3 = earlyWinner_3_1 ? beatsDO_1 : 3'h0; // @[Arbiter.scala 111:73]
  wire [8:0] _GEN_17 = {{6'd0}, maskedBeats_1_3}; // @[Arbiter.scala 112:44]
  wire [8:0] initBeats_3 = maskedBeats_0_3 | _GEN_17; // @[Arbiter.scala 112:44]
  wire  _sink_ACancel_earlyValid_T_8 = state_3_0 & portsDIO_filtered__1_valid | state_3_1 & portsDIO_filtered_1_1_valid; // @[Mux.scala 27:73]
  wire  sink_ACancel_7_earlyValid = idle_3 ? _T_196 : _sink_ACancel_earlyValid_T_8; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_20 = auto_in_1_d_ready & sink_ACancel_7_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [8:0] _GEN_18 = {{8'd0}, _beatsLeft_T_20}; // @[Arbiter.scala 113:52]
  wire [8:0] _beatsLeft_T_22 = beatsLeft_3 - _GEN_18; // @[Arbiter.scala 113:52]
  wire [63:0] _T_213 = muxStateEarly_3_0 ? auto_out_0_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_214 = muxStateEarly_3_1 ? auto_out_1_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_225 = muxStateEarly_3_0 ? auto_out_0_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_226 = muxStateEarly_3_1 ? out_2_1_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_231 = muxStateEarly_3_0 ? auto_out_0_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_232 = muxStateEarly_3_1 ? auto_out_1_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  reg [15:0] TLXbar_covState; // @[Register tracking TLXbar state]
  reg  TLXbar_covMap [0:65535]; // @[Coverage map for TLXbar]
  wire  TLXbar_covMap_read_en; // @[Coverage map for TLXbar]
  wire [15:0] TLXbar_covMap_read_addr; // @[Coverage map for TLXbar]
  wire  TLXbar_covMap_read_data; // @[Coverage map for TLXbar]
  wire  TLXbar_covMap_write_data; // @[Coverage map for TLXbar]
  wire [15:0] TLXbar_covMap_write_addr; // @[Coverage map for TLXbar]
  wire  TLXbar_covMap_write_mask; // @[Coverage map for TLXbar]
  wire  TLXbar_covMap_write_en; // @[Coverage map for TLXbar]
  reg [29:0] TLXbar_covSum; // @[Sum of coverage map]
  wire [1:0] readys_mask_shl;
  wire [15:0] readys_mask_pad;
  wire [2:0] state_3_1_shl;
  wire [15:0] state_3_1_pad;
  wire [4:0] readys_mask_1_shl;
  wire [15:0] readys_mask_1_pad;
  wire [6:0] readys_mask_2_shl;
  wire [15:0] readys_mask_2_pad;
  wire [7:0] state_1_0_shl;
  wire [15:0] state_1_0_pad;
  wire [8:0] state__0_shl;
  wire [15:0] state__0_pad;
  wire [9:0] state_3_0_shl;
  wire [15:0] state_3_0_pad;
  wire [10:0] state__1_shl;
  wire [15:0] state__1_pad;
  wire [11:0] state_1_1_shl;
  wire [15:0] state_1_1_pad;
  wire [12:0] state_2_0_shl;
  wire [15:0] state_2_0_pad;
  wire [14:0] readys_mask_3_shl;
  wire [15:0] readys_mask_3_pad;
  wire [15:0] state_2_1_shl;
  wire [15:0] state_2_1_pad;
  wire [15:0] TLXbar_xor8;
  wire [15:0] TLXbar_xor3;
  wire [15:0] TLXbar_xor10;
  wire [15:0] TLXbar_xor4;
  wire [15:0] TLXbar_xor1;
  wire [15:0] TLXbar_xor12;
  wire [15:0] TLXbar_xor5;
  wire [15:0] TLXbar_xor14;
  wire [15:0] TLXbar_xor6;
  wire [15:0] TLXbar_xor2;
  wire [15:0] TLXbar_xor0;
  assign auto_in_1_a_ready = requestAIO_1_0 & portsAOI_filtered_1_0_ready | requestAIO_1_1 & portsAOI_filtered_1_1_ready
    ; // @[Mux.scala 27:73]
  assign auto_in_1_d_valid = idle_3 ? _T_196 : _sink_ACancel_earlyValid_T_8; // @[Arbiter.scala 125:29]
  assign auto_in_1_d_bits_opcode = _T_231 | _T_232; // @[Mux.scala 27:73]
  assign auto_in_1_d_bits_size = _T_225 | _T_226; // @[Mux.scala 27:73]
  assign auto_in_1_d_bits_source = sink_ACancel_7_bits_source[5:0]; // @[Xbar.scala 228:69]
  assign auto_in_1_d_bits_denied = muxStateEarly_3_0 & auto_out_0_d_bits_denied | muxStateEarly_3_1 &
    auto_out_1_d_bits_denied; // @[Mux.scala 27:73]
  assign auto_in_1_d_bits_data = _T_213 | _T_214; // @[Mux.scala 27:73]
  assign auto_in_1_d_bits_corrupt = muxStateEarly_3_0 & auto_out_0_d_bits_corrupt | muxStateEarly_3_1 &
    auto_out_1_d_bits_corrupt; // @[Mux.scala 27:73]
  assign auto_in_0_a_ready = requestAIO_0_0 & portsAOI_filtered__0_ready | requestAIO_0_1 & portsAOI_filtered__1_ready; // @[Mux.scala 27:73]
  assign auto_in_0_d_valid = idle_2 ? _T_148 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_in_0_d_bits_opcode = _T_183 | _T_184; // @[Mux.scala 27:73]
  assign auto_in_0_d_bits_size = _T_177 | _T_178; // @[Mux.scala 27:73]
  assign auto_in_0_d_bits_source = sink_ACancel_5_bits_source[3:0]; // @[Xbar.scala 228:69]
  assign auto_in_0_d_bits_denied = muxStateEarly_2_0 & auto_out_0_d_bits_denied | muxStateEarly_2_1 &
    auto_out_1_d_bits_denied; // @[Mux.scala 27:73]
  assign auto_in_0_d_bits_data = _T_165 | _T_166; // @[Mux.scala 27:73]
  assign auto_in_0_d_bits_corrupt = muxStateEarly_2_0 & auto_out_0_d_bits_corrupt | muxStateEarly_2_1 &
    auto_out_1_d_bits_corrupt; // @[Mux.scala 27:73]
  assign auto_out_1_a_valid = idle_1 ? _T_79 : _out_1_a_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_out_1_a_bits_opcode = _T_135 | _T_136; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_size = out_2_1_a_bits_size[2:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_1_a_bits_source = _T_126 | _T_127; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_address = _T_123 | _T_124; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_user_amba_prot_bufferable = muxStateEarly_1_0 & auto_in_0_a_bits_user_amba_prot_bufferable |
    muxStateEarly_1_1 & auto_in_1_a_bits_user_amba_prot_bufferable; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_user_amba_prot_modifiable = muxStateEarly_1_0 & auto_in_0_a_bits_user_amba_prot_modifiable |
    muxStateEarly_1_1 & auto_in_1_a_bits_user_amba_prot_modifiable; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_user_amba_prot_readalloc = muxStateEarly_1_0 & auto_in_0_a_bits_user_amba_prot_readalloc |
    muxStateEarly_1_1 & auto_in_1_a_bits_user_amba_prot_readalloc; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_user_amba_prot_writealloc = muxStateEarly_1_0 & auto_in_0_a_bits_user_amba_prot_writealloc |
    muxStateEarly_1_1 & auto_in_1_a_bits_user_amba_prot_writealloc; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_user_amba_prot_privileged = muxStateEarly_1_0 & auto_in_0_a_bits_user_amba_prot_privileged |
    muxStateEarly_1_1 & auto_in_1_a_bits_user_amba_prot_privileged; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_user_amba_prot_secure = muxStateEarly_1_0 & auto_in_0_a_bits_user_amba_prot_secure |
    muxStateEarly_1_1 & auto_in_1_a_bits_user_amba_prot_secure; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_user_amba_prot_fetch = muxStateEarly_1_0 & auto_in_0_a_bits_user_amba_prot_fetch |
    muxStateEarly_1_1 & auto_in_1_a_bits_user_amba_prot_fetch; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_mask = _T_99 | _T_100; // @[Mux.scala 27:73]
  assign auto_out_1_a_bits_data = _T_96 | _T_97; // @[Mux.scala 27:73]
  assign auto_out_1_d_ready = requestDOI_1_0 & out_9_ready | requestDOI_1_1 & out_13_ready; // @[Mux.scala 27:73]
  assign auto_out_0_a_valid = idle ? _T_10 : _out_0_a_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_out_0_a_bits_opcode = _T_66 | _T_67; // @[Mux.scala 27:73]
  assign auto_out_0_a_bits_param = _T_63 | _T_64; // @[Mux.scala 27:73]
  assign auto_out_0_a_bits_size = _T_60 | _T_61; // @[Mux.scala 27:73]
  assign auto_out_0_a_bits_source = _T_57 | _T_58; // @[Mux.scala 27:73]
  assign auto_out_0_a_bits_address = out_2_0_a_bits_address[30:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_0_a_bits_mask = _T_30 | _T_31; // @[Mux.scala 27:73]
  assign auto_out_0_a_bits_data = _T_27 | _T_28; // @[Mux.scala 27:73]
  assign auto_out_0_d_ready = requestDOI_0_0 & out_8_ready | requestDOI_0_1 & out_12_ready; // @[Mux.scala 27:73]
  assign TLXbar_covMap_read_en = 1'h1;
  assign TLXbar_covMap_read_addr = TLXbar_covState;
  assign TLXbar_covMap_read_data = TLXbar_covMap[TLXbar_covMap_read_addr]; // @[Coverage map for TLXbar]
  assign TLXbar_covMap_write_data = 1'h1;
  assign TLXbar_covMap_write_addr = TLXbar_covState;
  assign TLXbar_covMap_write_mask = 1'h1;
  assign TLXbar_covMap_write_en = ~metaReset;
  assign readys_mask_shl = readys_mask;
  assign readys_mask_pad = {14'h0,readys_mask_shl};
  assign state_3_1_shl = {state_3_1, 2'h0};
  assign state_3_1_pad = {13'h0,state_3_1_shl};
  assign readys_mask_1_shl = {readys_mask_1, 3'h0};
  assign readys_mask_1_pad = {11'h0,readys_mask_1_shl};
  assign readys_mask_2_shl = {readys_mask_2, 5'h0};
  assign readys_mask_2_pad = {9'h0,readys_mask_2_shl};
  assign state_1_0_shl = {state_1_0, 7'h0};
  assign state_1_0_pad = {8'h0,state_1_0_shl};
  assign state__0_shl = {state__0, 8'h0};
  assign state__0_pad = {7'h0,state__0_shl};
  assign state_3_0_shl = {state_3_0, 9'h0};
  assign state_3_0_pad = {6'h0,state_3_0_shl};
  assign state__1_shl = {state__1, 10'h0};
  assign state__1_pad = {5'h0,state__1_shl};
  assign state_1_1_shl = {state_1_1, 11'h0};
  assign state_1_1_pad = {4'h0,state_1_1_shl};
  assign state_2_0_shl = {state_2_0, 12'h0};
  assign state_2_0_pad = {3'h0,state_2_0_shl};
  assign readys_mask_3_shl = {readys_mask_3, 13'h0};
  assign readys_mask_3_pad = {1'h0,readys_mask_3_shl};
  assign state_2_1_shl = {state_2_1, 15'h0};
  assign state_2_1_pad = state_2_1_shl;
  assign TLXbar_xor8 = state_3_1_pad ^ readys_mask_1_pad;
  assign TLXbar_xor3 = readys_mask_pad ^ TLXbar_xor8;
  assign TLXbar_xor10 = state_1_0_pad ^ state__0_pad;
  assign TLXbar_xor4 = readys_mask_2_pad ^ TLXbar_xor10;
  assign TLXbar_xor1 = TLXbar_xor3 ^ TLXbar_xor4;
  assign TLXbar_xor12 = state__1_pad ^ state_1_1_pad;
  assign TLXbar_xor5 = state_3_0_pad ^ TLXbar_xor12;
  assign TLXbar_xor14 = readys_mask_3_pad ^ state_2_1_pad;
  assign TLXbar_xor6 = state_2_0_pad ^ TLXbar_xor14;
  assign TLXbar_xor2 = TLXbar_xor5 ^ TLXbar_xor6;
  assign TLXbar_xor0 = TLXbar_xor1 ^ TLXbar_xor2;
  assign io_covSum = TLXbar_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft_2 <= 9'h0; // @[Arbiter.scala 87:30]
    end else if (latch_2) begin
      beatsLeft_2 <= initBeats_2;
    end else begin
      beatsLeft_2 <= _beatsLeft_T_16;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask_2 <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (latch_2 & |readys_valid_2) begin
      readys_mask_2 <= _readys_mask_T_13;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_2_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_2) begin
      state_2_0 <= earlyWinner_2_0;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_2_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_2) begin
      state_2_1 <= earlyWinner_2_1;
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft_3 <= 9'h0; // @[Arbiter.scala 87:30]
    end else if (latch_3) begin
      beatsLeft_3 <= initBeats_3;
    end else begin
      beatsLeft_3 <= _beatsLeft_T_22;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask_3 <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (latch_3 & |readys_valid_3) begin
      readys_mask_3 <= _readys_mask_T_18;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_3_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_3) begin
      state_3_0 <= earlyWinner_3_0;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_3_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_3) begin
      state_3_1 <= earlyWinner_3_1;
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 9'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin
      beatsLeft <= initBeats;
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (latch & |readys_valid) begin
      readys_mask <= _readys_mask_T_3;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state__0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state__0 <= earlyWinner__0;
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft_1 <= 9'h0; // @[Arbiter.scala 87:30]
    end else if (latch_1) begin
      beatsLeft_1 <= initBeats_1;
    end else begin
      beatsLeft_1 <= _beatsLeft_T_10;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask_1 <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (latch_1 & |readys_valid_1) begin
      readys_mask_1 <= _readys_mask_T_8;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin
      state_1_0 <= earlyWinner_1_0;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state__1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state__1 <= earlyWinner__1;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin
      state_1_1 <= earlyWinner_1_1;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Arbiter.scala 22:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner__0 | ~earlyWinner__1) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~earlyWinner__0 | ~earlyWinner__1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(portsAOI_filtered__0_earlyValid | portsAOI_filtered_1_0_earlyValid) | (earlyWinner__0 | earlyWinner__1))
           & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~(portsAOI_filtered__0_earlyValid | portsAOI_filtered_1_0_earlyValid) | (earlyWinner__0 |
          earlyWinner__1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_11 | _T_10) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(_T_11 | _T_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Arbiter.scala 22:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_1_0 | ~earlyWinner_1_1) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~earlyWinner_1_0 | ~earlyWinner_1_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(portsAOI_filtered__1_earlyValid | portsAOI_filtered_1_1_earlyValid) | (earlyWinner_1_0 | earlyWinner_1_1
          )) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~(portsAOI_filtered__1_earlyValid | portsAOI_filtered_1_1_earlyValid) | (earlyWinner_1_0 |
          earlyWinner_1_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_80 | _T_79) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(_T_80 | _T_79)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Arbiter.scala 22:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_2_0 | ~earlyWinner_2_1) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~earlyWinner_2_0 | ~earlyWinner_2_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(portsDIO_filtered__0_valid | portsDIO_filtered_1_0_valid) | (earlyWinner_2_0 | earlyWinner_2_1)) &
          _readys_T_3) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~(portsDIO_filtered__0_valid | portsDIO_filtered_1_0_valid) | (earlyWinner_2_0 |
          earlyWinner_2_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_149 | _T_148) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(_T_149 | _T_148)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Arbiter.scala 22:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_3_0 | ~earlyWinner_3_1) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~earlyWinner_3_0 | ~earlyWinner_3_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(portsDIO_filtered__1_valid | portsDIO_filtered_1_1_valid) | (earlyWinner_3_0 | earlyWinner_3_1)) &
          _readys_T_3) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~(portsDIO_filtered__1_valid | portsDIO_filtered_1_1_valid) | (earlyWinner_3_0 |
          earlyWinner_3_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_197 | _T_196) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(_T_197 | _T_196)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    TLXbar_covState <= TLXbar_xor0;
    if (TLXbar_covMap_write_en & TLXbar_covMap_write_mask) begin
      TLXbar_covMap[TLXbar_covMap_write_addr] <= TLXbar_covMap_write_data; // @[Coverage map for TLXbar]
    end
    if (!(TLXbar_covMap_read_data | metaReset)) begin
      TLXbar_covSum <= TLXbar_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 65536; initvar = initvar+1)
    TLXbar_covMap[initvar] = 0; //_17[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft_2 = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  readys_mask_2 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  state_2_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_2_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  beatsLeft_3 = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  readys_mask_3 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  state_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  beatsLeft = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  readys_mask = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  state__0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  beatsLeft_1 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  readys_mask_1 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  state_1_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state__1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_1_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  TLXbar_covState = 0; //_16[15:0];
  _RAND_18 = {1{`RANDOM}};
  TLXbar_covSum = 0; //_18[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFIFOFixer(
  output        auto_in_1_a_ready,
  input         auto_in_1_a_valid,
  input  [2:0]  auto_in_1_a_bits_opcode,
  input  [2:0]  auto_in_1_a_bits_param,
  input  [3:0]  auto_in_1_a_bits_size,
  input  [5:0]  auto_in_1_a_bits_source,
  input  [31:0] auto_in_1_a_bits_address,
  input         auto_in_1_a_bits_user_amba_prot_bufferable,
  input         auto_in_1_a_bits_user_amba_prot_modifiable,
  input         auto_in_1_a_bits_user_amba_prot_readalloc,
  input         auto_in_1_a_bits_user_amba_prot_writealloc,
  input         auto_in_1_a_bits_user_amba_prot_privileged,
  input         auto_in_1_a_bits_user_amba_prot_secure,
  input         auto_in_1_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_1_a_bits_mask,
  input  [63:0] auto_in_1_a_bits_data,
  input         auto_in_1_d_ready,
  output        auto_in_1_d_valid,
  output [2:0]  auto_in_1_d_bits_opcode,
  output [3:0]  auto_in_1_d_bits_size,
  output [5:0]  auto_in_1_d_bits_source,
  output        auto_in_1_d_bits_denied,
  output [63:0] auto_in_1_d_bits_data,
  output        auto_in_1_d_bits_corrupt,
  output        auto_in_0_a_ready,
  input         auto_in_0_a_valid,
  input  [2:0]  auto_in_0_a_bits_opcode,
  input  [2:0]  auto_in_0_a_bits_param,
  input  [3:0]  auto_in_0_a_bits_size,
  input  [3:0]  auto_in_0_a_bits_source,
  input  [31:0] auto_in_0_a_bits_address,
  input         auto_in_0_a_bits_user_amba_prot_bufferable,
  input         auto_in_0_a_bits_user_amba_prot_modifiable,
  input         auto_in_0_a_bits_user_amba_prot_readalloc,
  input         auto_in_0_a_bits_user_amba_prot_writealloc,
  input         auto_in_0_a_bits_user_amba_prot_privileged,
  input         auto_in_0_a_bits_user_amba_prot_secure,
  input         auto_in_0_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_0_a_bits_mask,
  input  [63:0] auto_in_0_a_bits_data,
  input         auto_in_0_d_ready,
  output        auto_in_0_d_valid,
  output [2:0]  auto_in_0_d_bits_opcode,
  output [3:0]  auto_in_0_d_bits_size,
  output [3:0]  auto_in_0_d_bits_source,
  output        auto_in_0_d_bits_denied,
  output [63:0] auto_in_0_d_bits_data,
  output        auto_in_0_d_bits_corrupt,
  input         auto_out_1_a_ready,
  output        auto_out_1_a_valid,
  output [2:0]  auto_out_1_a_bits_opcode,
  output [2:0]  auto_out_1_a_bits_param,
  output [3:0]  auto_out_1_a_bits_size,
  output [5:0]  auto_out_1_a_bits_source,
  output [31:0] auto_out_1_a_bits_address,
  output        auto_out_1_a_bits_user_amba_prot_bufferable,
  output        auto_out_1_a_bits_user_amba_prot_modifiable,
  output        auto_out_1_a_bits_user_amba_prot_readalloc,
  output        auto_out_1_a_bits_user_amba_prot_writealloc,
  output        auto_out_1_a_bits_user_amba_prot_privileged,
  output        auto_out_1_a_bits_user_amba_prot_secure,
  output        auto_out_1_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_1_a_bits_mask,
  output [63:0] auto_out_1_a_bits_data,
  output        auto_out_1_d_ready,
  input         auto_out_1_d_valid,
  input  [2:0]  auto_out_1_d_bits_opcode,
  input  [3:0]  auto_out_1_d_bits_size,
  input  [5:0]  auto_out_1_d_bits_source,
  input         auto_out_1_d_bits_denied,
  input  [63:0] auto_out_1_d_bits_data,
  input         auto_out_1_d_bits_corrupt,
  input         auto_out_0_a_ready,
  output        auto_out_0_a_valid,
  output [2:0]  auto_out_0_a_bits_opcode,
  output [2:0]  auto_out_0_a_bits_param,
  output [3:0]  auto_out_0_a_bits_size,
  output [3:0]  auto_out_0_a_bits_source,
  output [31:0] auto_out_0_a_bits_address,
  output        auto_out_0_a_bits_user_amba_prot_bufferable,
  output        auto_out_0_a_bits_user_amba_prot_modifiable,
  output        auto_out_0_a_bits_user_amba_prot_readalloc,
  output        auto_out_0_a_bits_user_amba_prot_writealloc,
  output        auto_out_0_a_bits_user_amba_prot_privileged,
  output        auto_out_0_a_bits_user_amba_prot_secure,
  output        auto_out_0_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_0_a_bits_mask,
  output [63:0] auto_out_0_a_bits_data,
  output        auto_out_0_d_ready,
  input         auto_out_0_d_valid,
  input  [2:0]  auto_out_0_d_bits_opcode,
  input  [3:0]  auto_out_0_d_bits_size,
  input  [3:0]  auto_out_0_d_bits_source,
  input         auto_out_0_d_bits_denied,
  input  [63:0] auto_out_0_d_bits_data,
  input         auto_out_0_d_bits_corrupt,
  output [29:0] io_covSum
);
  wire [29:0] TLFIFOFixer_covSum;
  assign auto_in_1_a_ready = auto_out_1_a_ready; // @[FIFOFixer.scala 88:33]
  assign auto_in_1_d_valid = auto_out_1_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_opcode = auto_out_1_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_size = auto_out_1_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_source = auto_out_1_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_denied = auto_out_1_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_data = auto_out_1_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_1_d_bits_corrupt = auto_out_1_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_0_a_ready = auto_out_0_a_ready; // @[FIFOFixer.scala 88:33]
  assign auto_in_0_d_valid = auto_out_0_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_0_d_bits_opcode = auto_out_0_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_0_d_bits_size = auto_out_0_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_0_d_bits_source = auto_out_0_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_0_d_bits_denied = auto_out_0_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_0_d_bits_data = auto_out_0_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_0_d_bits_corrupt = auto_out_0_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_1_a_valid = auto_in_1_a_valid; // @[FIFOFixer.scala 87:33]
  assign auto_out_1_a_bits_opcode = auto_in_1_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_param = auto_in_1_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_size = auto_in_1_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_source = auto_in_1_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_address = auto_in_1_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_user_amba_prot_bufferable = auto_in_1_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_user_amba_prot_modifiable = auto_in_1_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_user_amba_prot_readalloc = auto_in_1_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_user_amba_prot_writealloc = auto_in_1_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_user_amba_prot_privileged = auto_in_1_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_user_amba_prot_secure = auto_in_1_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_user_amba_prot_fetch = auto_in_1_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_mask = auto_in_1_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_data = auto_in_1_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_d_ready = auto_in_1_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_valid = auto_in_0_a_valid; // @[FIFOFixer.scala 87:33]
  assign auto_out_0_a_bits_opcode = auto_in_0_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_param = auto_in_0_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_size = auto_in_0_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_source = auto_in_0_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_address = auto_in_0_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_user_amba_prot_bufferable = auto_in_0_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_user_amba_prot_modifiable = auto_in_0_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_user_amba_prot_readalloc = auto_in_0_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_user_amba_prot_writealloc = auto_in_0_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_user_amba_prot_privileged = auto_in_0_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_user_amba_prot_secure = auto_in_0_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_user_amba_prot_fetch = auto_in_0_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_mask = auto_in_0_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_data = auto_in_0_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_d_ready = auto_in_0_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLFIFOFixer_covSum = 30'h0;
  assign io_covSum = TLFIFOFixer_covSum;
endmodule
module SystemBus(
  output        auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_ready,
  input         auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_valid,
  input  [2:0]  auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_opcode,
  input  [2:0]  auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_param,
  input  [3:0]  auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_size,
  input  [5:0]  auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_source,
  input  [31:0] auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_address,
  input         auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_bufferable,
  input         auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_modifiable,
  input         auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_readalloc,
  input         auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_writealloc,
  input         auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_privileged,
  input         auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_secure,
  input         auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_mask,
  input  [63:0] auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_data,
  input         auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_ready,
  output        auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_valid,
  output [2:0]  auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_opcode,
  output [3:0]  auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_size,
  output [5:0]  auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_source,
  output        auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_denied,
  output [63:0] auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_data,
  output        auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_corrupt,
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready,
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid,
  output [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode,
  output [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size,
  output [6:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source,
  output [31:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address,
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_bufferable,
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_modifiable,
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_readalloc,
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_writealloc,
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_privileged,
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_secure,
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask,
  output [63:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data,
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready,
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid,
  input  [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode,
  input  [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size,
  input  [6:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source,
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied,
  input  [63:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data,
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt,
  output        auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready,
  input         auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid,
  input  [2:0]  auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode,
  input  [2:0]  auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param,
  input  [3:0]  auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size,
  input  [3:0]  auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source,
  input  [31:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address,
  input         auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_bufferable,
  input         auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_modifiable,
  input         auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_readalloc,
  input         auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_writealloc,
  input         auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_privileged,
  input         auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_secure,
  input         auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask,
  input  [63:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data,
  input         auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready,
  output        auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid,
  output [2:0]  auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode,
  output [3:0]  auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size,
  output [3:0]  auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source,
  output        auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied,
  output [63:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data,
  output        auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt,
  input         auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready,
  output        auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid,
  output [2:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode,
  output [2:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param,
  output [3:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size,
  output [6:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source,
  output [30:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address,
  output [7:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask,
  output [63:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data,
  output        auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready,
  input         auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid,
  input  [2:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode,
  input  [3:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size,
  input  [6:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source,
  input         auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied,
  input  [63:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data,
  input         auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt,
  output        auto_fixedClockNode_out_1_clock,
  output        auto_fixedClockNode_out_1_reset,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock,
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset,
  output        auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock,
  output        auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset,
  output        auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock,
  output        auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset,
  output        auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock,
  output        auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset,
  output        auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock,
  output        auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset,
  output        auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock,
  output        auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_clock;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_reset;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_clock;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_reset;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_clock;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_reset;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_clock;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_reset;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_clock;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_reset;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_clock;
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_reset;
  wire  subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_clock;
  wire  subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_reset;
  wire  subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_clock;
  wire  subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_reset;
  wire  subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_clock;
  wire  subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_reset;
  wire  subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_clock;
  wire  subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_reset;
  wire  subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_clock;
  wire  subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_reset;
  wire  subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_clock;
  wire  subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_reset;
  wire  clockGroup_auto_in_member_subsystem_sbus_0_clock;
  wire  clockGroup_auto_in_member_subsystem_sbus_0_reset;
  wire  clockGroup_auto_out_clock;
  wire  clockGroup_auto_out_reset;
  wire  fixedClockNode_auto_in_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_in_reset; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_2_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_2_reset; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_1_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_1_reset; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_0_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_0_reset; // @[ClockGroup.scala 106:107]
  wire [29:0] fixedClockNode_io_covSum; // @[ClockGroup.scala 106:107]
  wire  system_bus_xbar_clock; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_reset; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_a_ready; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_a_valid; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_1_a_bits_opcode; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_1_a_bits_param; // @[SystemBus.scala 40:43]
  wire [3:0] system_bus_xbar_auto_in_1_a_bits_size; // @[SystemBus.scala 40:43]
  wire [5:0] system_bus_xbar_auto_in_1_a_bits_source; // @[SystemBus.scala 40:43]
  wire [31:0] system_bus_xbar_auto_in_1_a_bits_address; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_a_bits_user_amba_prot_bufferable; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_a_bits_user_amba_prot_modifiable; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_a_bits_user_amba_prot_readalloc; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_a_bits_user_amba_prot_writealloc; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_a_bits_user_amba_prot_privileged; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_a_bits_user_amba_prot_secure; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_a_bits_user_amba_prot_fetch; // @[SystemBus.scala 40:43]
  wire [7:0] system_bus_xbar_auto_in_1_a_bits_mask; // @[SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_in_1_a_bits_data; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_d_ready; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_d_valid; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_1_d_bits_opcode; // @[SystemBus.scala 40:43]
  wire [3:0] system_bus_xbar_auto_in_1_d_bits_size; // @[SystemBus.scala 40:43]
  wire [5:0] system_bus_xbar_auto_in_1_d_bits_source; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_d_bits_denied; // @[SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_in_1_d_bits_data; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_1_d_bits_corrupt; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_a_ready; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_a_valid; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_0_a_bits_opcode; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_0_a_bits_param; // @[SystemBus.scala 40:43]
  wire [3:0] system_bus_xbar_auto_in_0_a_bits_size; // @[SystemBus.scala 40:43]
  wire [3:0] system_bus_xbar_auto_in_0_a_bits_source; // @[SystemBus.scala 40:43]
  wire [31:0] system_bus_xbar_auto_in_0_a_bits_address; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_a_bits_user_amba_prot_bufferable; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_a_bits_user_amba_prot_modifiable; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_a_bits_user_amba_prot_readalloc; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_a_bits_user_amba_prot_writealloc; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_a_bits_user_amba_prot_privileged; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_a_bits_user_amba_prot_secure; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_a_bits_user_amba_prot_fetch; // @[SystemBus.scala 40:43]
  wire [7:0] system_bus_xbar_auto_in_0_a_bits_mask; // @[SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_in_0_a_bits_data; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_d_ready; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_d_valid; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_0_d_bits_opcode; // @[SystemBus.scala 40:43]
  wire [3:0] system_bus_xbar_auto_in_0_d_bits_size; // @[SystemBus.scala 40:43]
  wire [3:0] system_bus_xbar_auto_in_0_d_bits_source; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_d_bits_denied; // @[SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_in_0_d_bits_data; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_0_d_bits_corrupt; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_ready; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_valid; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_a_bits_opcode; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_a_bits_size; // @[SystemBus.scala 40:43]
  wire [6:0] system_bus_xbar_auto_out_1_a_bits_source; // @[SystemBus.scala 40:43]
  wire [31:0] system_bus_xbar_auto_out_1_a_bits_address; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_bits_user_amba_prot_bufferable; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_bits_user_amba_prot_modifiable; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_bits_user_amba_prot_readalloc; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_bits_user_amba_prot_writealloc; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_bits_user_amba_prot_privileged; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_bits_user_amba_prot_secure; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_bits_user_amba_prot_fetch; // @[SystemBus.scala 40:43]
  wire [7:0] system_bus_xbar_auto_out_1_a_bits_mask; // @[SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_out_1_a_bits_data; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_d_ready; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_d_valid; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_d_bits_opcode; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_d_bits_size; // @[SystemBus.scala 40:43]
  wire [6:0] system_bus_xbar_auto_out_1_d_bits_source; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_d_bits_denied; // @[SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_out_1_d_bits_data; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_d_bits_corrupt; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_a_ready; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_a_valid; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_0_a_bits_opcode; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_0_a_bits_param; // @[SystemBus.scala 40:43]
  wire [3:0] system_bus_xbar_auto_out_0_a_bits_size; // @[SystemBus.scala 40:43]
  wire [6:0] system_bus_xbar_auto_out_0_a_bits_source; // @[SystemBus.scala 40:43]
  wire [30:0] system_bus_xbar_auto_out_0_a_bits_address; // @[SystemBus.scala 40:43]
  wire [7:0] system_bus_xbar_auto_out_0_a_bits_mask; // @[SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_out_0_a_bits_data; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_d_ready; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_d_valid; // @[SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_0_d_bits_opcode; // @[SystemBus.scala 40:43]
  wire [3:0] system_bus_xbar_auto_out_0_d_bits_size; // @[SystemBus.scala 40:43]
  wire [6:0] system_bus_xbar_auto_out_0_d_bits_source; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_d_bits_denied; // @[SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_out_0_d_bits_data; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_d_bits_corrupt; // @[SystemBus.scala 40:43]
  wire [29:0] system_bus_xbar_io_covSum; // @[SystemBus.scala 40:43]
  wire  system_bus_xbar_metaReset; // @[SystemBus.scala 40:43]
  wire  fixer_auto_in_1_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_1_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_1_a_bits_param; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_1_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_in_1_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_in_1_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_in_1_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_1_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_1_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_1_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_in_1_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_1_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_1_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_0_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_0_a_bits_param; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_0_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_0_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_in_0_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_in_0_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_0_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_0_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_0_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_0_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_0_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_0_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_1_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_1_a_bits_param; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_1_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_out_1_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_out_1_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_out_1_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_1_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_1_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_1_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_out_1_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_1_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_1_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_0_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_0_a_bits_param; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_0_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_0_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_out_0_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_out_0_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_0_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_0_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_0_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_0_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_0_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_0_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire [29:0] fixer_io_covSum; // @[FIFOFixer.scala 144:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_ready;
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_param;
  wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_source;
  wire [30:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_address;
  wire [7:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_data;
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_ready;
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_opcode;
  wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_source;
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_data;
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_ready;
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_param;
  wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_source;
  wire [30:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_address;
  wire [7:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_data;
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_ready;
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_opcode;
  wire [3:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_source;
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_data;
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_ready;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_param;
  wire [3:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_source;
  wire [30:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_address;
  wire [7:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_data;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_ready;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_opcode;
  wire [3:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_source;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_data;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_ready;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_param;
  wire [3:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_source;
  wire [30:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_address;
  wire [7:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_data;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_ready;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_opcode;
  wire [3:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_source;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_data;
  wire  coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_corrupt;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_ready;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_valid;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_opcode;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_param;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_size;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_source;
  wire [31:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_address;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_bufferable;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_modifiable;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_readalloc;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_writealloc;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_privileged;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_secure;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_mask;
  wire [63:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_data;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_ready;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_valid;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_opcode;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_size;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_source;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_denied;
  wire [63:0] coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_data;
  wire  coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_corrupt;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_ready;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_valid;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_opcode;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_param;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_size;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_source;
  wire [31:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_address;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_bufferable;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_modifiable;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_readalloc;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_writealloc;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_privileged;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_secure;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_mask;
  wire [63:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_data;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_ready;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_valid;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_opcode;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_size;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_source;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_denied;
  wire [63:0] coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_data;
  wire  coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_corrupt;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_ready;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_valid;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_opcode;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_param;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_size;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_source;
  wire [31:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_address;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_bufferable;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_modifiable;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_readalloc;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_writealloc;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_privileged;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_secure;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_mask;
  wire [63:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_data;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_ready;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_valid;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_opcode;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_size;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_source;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_denied;
  wire [63:0] coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_data;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_corrupt;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_ready;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_valid;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_opcode;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_param;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_size;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_source;
  wire [31:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_address;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_bufferable;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_modifiable;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_readalloc;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_writealloc;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_privileged;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_secure;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_mask;
  wire [63:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_data;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_ready;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_valid;
  wire [2:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_opcode;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_size;
  wire [3:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_source;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_denied;
  wire [63:0] coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_data;
  wire  coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_ready;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_source;
  wire [31:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_address;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_bufferable;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_modifiable;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_readalloc;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_writealloc;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_privileged;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_secure;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_data;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_d_ready;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_source;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_data;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_ready;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_source;
  wire [31:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_address;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_bufferable;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_modifiable;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_readalloc;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_writealloc;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_privileged;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_secure;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_data;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_d_ready;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_source;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_data;
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_a_ready;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_source;
  wire [31:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_address;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_bufferable;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_modifiable;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_readalloc;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_writealloc;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_privileged;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_secure;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_data;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_d_ready;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_source;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_data;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_a_ready;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_source;
  wire [31:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_address;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_bufferable;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_modifiable;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_readalloc;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_writealloc;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_privileged;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_secure;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_data;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_d_ready;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_source;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_data;
  wire  coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_corrupt;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_ready;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_valid;
  wire [2:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_opcode;
  wire [2:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_param;
  wire [3:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_size;
  wire [5:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_source;
  wire [31:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_address;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_bufferable;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_modifiable;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_readalloc;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_writealloc;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_privileged;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_secure;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_mask;
  wire [63:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_data;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_ready;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_valid;
  wire [2:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_opcode;
  wire [3:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_size;
  wire [5:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_source;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_denied;
  wire [63:0] coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_data;
  wire  coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_corrupt;
  wire  coupler_from_cva6_tile_auto_tl_out_a_ready;
  wire  coupler_from_cva6_tile_auto_tl_out_a_valid;
  wire [2:0] coupler_from_cva6_tile_auto_tl_out_a_bits_opcode;
  wire [2:0] coupler_from_cva6_tile_auto_tl_out_a_bits_param;
  wire [3:0] coupler_from_cva6_tile_auto_tl_out_a_bits_size;
  wire [5:0] coupler_from_cva6_tile_auto_tl_out_a_bits_source;
  wire [31:0] coupler_from_cva6_tile_auto_tl_out_a_bits_address;
  wire  coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_bufferable;
  wire  coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_modifiable;
  wire  coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_readalloc;
  wire  coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_writealloc;
  wire  coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_privileged;
  wire  coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_secure;
  wire  coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_from_cva6_tile_auto_tl_out_a_bits_mask;
  wire [63:0] coupler_from_cva6_tile_auto_tl_out_a_bits_data;
  wire  coupler_from_cva6_tile_auto_tl_out_d_ready;
  wire  coupler_from_cva6_tile_auto_tl_out_d_valid;
  wire [2:0] coupler_from_cva6_tile_auto_tl_out_d_bits_opcode;
  wire [3:0] coupler_from_cva6_tile_auto_tl_out_d_bits_size;
  wire [5:0] coupler_from_cva6_tile_auto_tl_out_d_bits_source;
  wire  coupler_from_cva6_tile_auto_tl_out_d_bits_denied;
  wire [63:0] coupler_from_cva6_tile_auto_tl_out_d_bits_data;
  wire  coupler_from_cva6_tile_auto_tl_out_d_bits_corrupt;
  wire [29:0] SystemBus_covSum;
  wire [29:0] fixedClockNode_sum;
  wire [29:0] system_bus_xbar_sum;
  wire [29:0] fixer_sum;
  FixedClockBroadcast fixedClockNode ( // @[ClockGroup.scala 106:107]
    .auto_in_clock(fixedClockNode_auto_in_clock),
    .auto_in_reset(fixedClockNode_auto_in_reset),
    .auto_out_2_clock(fixedClockNode_auto_out_2_clock),
    .auto_out_2_reset(fixedClockNode_auto_out_2_reset),
    .auto_out_1_clock(fixedClockNode_auto_out_1_clock),
    .auto_out_1_reset(fixedClockNode_auto_out_1_reset),
    .auto_out_0_clock(fixedClockNode_auto_out_0_clock),
    .auto_out_0_reset(fixedClockNode_auto_out_0_reset),
    .io_covSum(fixedClockNode_io_covSum)
  );
  TLXbar system_bus_xbar ( // @[SystemBus.scala 40:43]
    .clock(system_bus_xbar_clock),
    .reset(system_bus_xbar_reset),
    .auto_in_1_a_ready(system_bus_xbar_auto_in_1_a_ready),
    .auto_in_1_a_valid(system_bus_xbar_auto_in_1_a_valid),
    .auto_in_1_a_bits_opcode(system_bus_xbar_auto_in_1_a_bits_opcode),
    .auto_in_1_a_bits_param(system_bus_xbar_auto_in_1_a_bits_param),
    .auto_in_1_a_bits_size(system_bus_xbar_auto_in_1_a_bits_size),
    .auto_in_1_a_bits_source(system_bus_xbar_auto_in_1_a_bits_source),
    .auto_in_1_a_bits_address(system_bus_xbar_auto_in_1_a_bits_address),
    .auto_in_1_a_bits_user_amba_prot_bufferable(system_bus_xbar_auto_in_1_a_bits_user_amba_prot_bufferable),
    .auto_in_1_a_bits_user_amba_prot_modifiable(system_bus_xbar_auto_in_1_a_bits_user_amba_prot_modifiable),
    .auto_in_1_a_bits_user_amba_prot_readalloc(system_bus_xbar_auto_in_1_a_bits_user_amba_prot_readalloc),
    .auto_in_1_a_bits_user_amba_prot_writealloc(system_bus_xbar_auto_in_1_a_bits_user_amba_prot_writealloc),
    .auto_in_1_a_bits_user_amba_prot_privileged(system_bus_xbar_auto_in_1_a_bits_user_amba_prot_privileged),
    .auto_in_1_a_bits_user_amba_prot_secure(system_bus_xbar_auto_in_1_a_bits_user_amba_prot_secure),
    .auto_in_1_a_bits_user_amba_prot_fetch(system_bus_xbar_auto_in_1_a_bits_user_amba_prot_fetch),
    .auto_in_1_a_bits_mask(system_bus_xbar_auto_in_1_a_bits_mask),
    .auto_in_1_a_bits_data(system_bus_xbar_auto_in_1_a_bits_data),
    .auto_in_1_d_ready(system_bus_xbar_auto_in_1_d_ready),
    .auto_in_1_d_valid(system_bus_xbar_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(system_bus_xbar_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_size(system_bus_xbar_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_source(system_bus_xbar_auto_in_1_d_bits_source),
    .auto_in_1_d_bits_denied(system_bus_xbar_auto_in_1_d_bits_denied),
    .auto_in_1_d_bits_data(system_bus_xbar_auto_in_1_d_bits_data),
    .auto_in_1_d_bits_corrupt(system_bus_xbar_auto_in_1_d_bits_corrupt),
    .auto_in_0_a_ready(system_bus_xbar_auto_in_0_a_ready),
    .auto_in_0_a_valid(system_bus_xbar_auto_in_0_a_valid),
    .auto_in_0_a_bits_opcode(system_bus_xbar_auto_in_0_a_bits_opcode),
    .auto_in_0_a_bits_param(system_bus_xbar_auto_in_0_a_bits_param),
    .auto_in_0_a_bits_size(system_bus_xbar_auto_in_0_a_bits_size),
    .auto_in_0_a_bits_source(system_bus_xbar_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(system_bus_xbar_auto_in_0_a_bits_address),
    .auto_in_0_a_bits_user_amba_prot_bufferable(system_bus_xbar_auto_in_0_a_bits_user_amba_prot_bufferable),
    .auto_in_0_a_bits_user_amba_prot_modifiable(system_bus_xbar_auto_in_0_a_bits_user_amba_prot_modifiable),
    .auto_in_0_a_bits_user_amba_prot_readalloc(system_bus_xbar_auto_in_0_a_bits_user_amba_prot_readalloc),
    .auto_in_0_a_bits_user_amba_prot_writealloc(system_bus_xbar_auto_in_0_a_bits_user_amba_prot_writealloc),
    .auto_in_0_a_bits_user_amba_prot_privileged(system_bus_xbar_auto_in_0_a_bits_user_amba_prot_privileged),
    .auto_in_0_a_bits_user_amba_prot_secure(system_bus_xbar_auto_in_0_a_bits_user_amba_prot_secure),
    .auto_in_0_a_bits_user_amba_prot_fetch(system_bus_xbar_auto_in_0_a_bits_user_amba_prot_fetch),
    .auto_in_0_a_bits_mask(system_bus_xbar_auto_in_0_a_bits_mask),
    .auto_in_0_a_bits_data(system_bus_xbar_auto_in_0_a_bits_data),
    .auto_in_0_d_ready(system_bus_xbar_auto_in_0_d_ready),
    .auto_in_0_d_valid(system_bus_xbar_auto_in_0_d_valid),
    .auto_in_0_d_bits_opcode(system_bus_xbar_auto_in_0_d_bits_opcode),
    .auto_in_0_d_bits_size(system_bus_xbar_auto_in_0_d_bits_size),
    .auto_in_0_d_bits_source(system_bus_xbar_auto_in_0_d_bits_source),
    .auto_in_0_d_bits_denied(system_bus_xbar_auto_in_0_d_bits_denied),
    .auto_in_0_d_bits_data(system_bus_xbar_auto_in_0_d_bits_data),
    .auto_in_0_d_bits_corrupt(system_bus_xbar_auto_in_0_d_bits_corrupt),
    .auto_out_1_a_ready(system_bus_xbar_auto_out_1_a_ready),
    .auto_out_1_a_valid(system_bus_xbar_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(system_bus_xbar_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_size(system_bus_xbar_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(system_bus_xbar_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(system_bus_xbar_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_user_amba_prot_bufferable(system_bus_xbar_auto_out_1_a_bits_user_amba_prot_bufferable),
    .auto_out_1_a_bits_user_amba_prot_modifiable(system_bus_xbar_auto_out_1_a_bits_user_amba_prot_modifiable),
    .auto_out_1_a_bits_user_amba_prot_readalloc(system_bus_xbar_auto_out_1_a_bits_user_amba_prot_readalloc),
    .auto_out_1_a_bits_user_amba_prot_writealloc(system_bus_xbar_auto_out_1_a_bits_user_amba_prot_writealloc),
    .auto_out_1_a_bits_user_amba_prot_privileged(system_bus_xbar_auto_out_1_a_bits_user_amba_prot_privileged),
    .auto_out_1_a_bits_user_amba_prot_secure(system_bus_xbar_auto_out_1_a_bits_user_amba_prot_secure),
    .auto_out_1_a_bits_user_amba_prot_fetch(system_bus_xbar_auto_out_1_a_bits_user_amba_prot_fetch),
    .auto_out_1_a_bits_mask(system_bus_xbar_auto_out_1_a_bits_mask),
    .auto_out_1_a_bits_data(system_bus_xbar_auto_out_1_a_bits_data),
    .auto_out_1_d_ready(system_bus_xbar_auto_out_1_d_ready),
    .auto_out_1_d_valid(system_bus_xbar_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(system_bus_xbar_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_size(system_bus_xbar_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(system_bus_xbar_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_denied(system_bus_xbar_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_data(system_bus_xbar_auto_out_1_d_bits_data),
    .auto_out_1_d_bits_corrupt(system_bus_xbar_auto_out_1_d_bits_corrupt),
    .auto_out_0_a_ready(system_bus_xbar_auto_out_0_a_ready),
    .auto_out_0_a_valid(system_bus_xbar_auto_out_0_a_valid),
    .auto_out_0_a_bits_opcode(system_bus_xbar_auto_out_0_a_bits_opcode),
    .auto_out_0_a_bits_param(system_bus_xbar_auto_out_0_a_bits_param),
    .auto_out_0_a_bits_size(system_bus_xbar_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(system_bus_xbar_auto_out_0_a_bits_source),
    .auto_out_0_a_bits_address(system_bus_xbar_auto_out_0_a_bits_address),
    .auto_out_0_a_bits_mask(system_bus_xbar_auto_out_0_a_bits_mask),
    .auto_out_0_a_bits_data(system_bus_xbar_auto_out_0_a_bits_data),
    .auto_out_0_d_ready(system_bus_xbar_auto_out_0_d_ready),
    .auto_out_0_d_valid(system_bus_xbar_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(system_bus_xbar_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_size(system_bus_xbar_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(system_bus_xbar_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_denied(system_bus_xbar_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_data(system_bus_xbar_auto_out_0_d_bits_data),
    .auto_out_0_d_bits_corrupt(system_bus_xbar_auto_out_0_d_bits_corrupt),
    .io_covSum(system_bus_xbar_io_covSum),
    .metaReset(system_bus_xbar_metaReset)
  );
  TLFIFOFixer fixer ( // @[FIFOFixer.scala 144:27]
    .auto_in_1_a_ready(fixer_auto_in_1_a_ready),
    .auto_in_1_a_valid(fixer_auto_in_1_a_valid),
    .auto_in_1_a_bits_opcode(fixer_auto_in_1_a_bits_opcode),
    .auto_in_1_a_bits_param(fixer_auto_in_1_a_bits_param),
    .auto_in_1_a_bits_size(fixer_auto_in_1_a_bits_size),
    .auto_in_1_a_bits_source(fixer_auto_in_1_a_bits_source),
    .auto_in_1_a_bits_address(fixer_auto_in_1_a_bits_address),
    .auto_in_1_a_bits_user_amba_prot_bufferable(fixer_auto_in_1_a_bits_user_amba_prot_bufferable),
    .auto_in_1_a_bits_user_amba_prot_modifiable(fixer_auto_in_1_a_bits_user_amba_prot_modifiable),
    .auto_in_1_a_bits_user_amba_prot_readalloc(fixer_auto_in_1_a_bits_user_amba_prot_readalloc),
    .auto_in_1_a_bits_user_amba_prot_writealloc(fixer_auto_in_1_a_bits_user_amba_prot_writealloc),
    .auto_in_1_a_bits_user_amba_prot_privileged(fixer_auto_in_1_a_bits_user_amba_prot_privileged),
    .auto_in_1_a_bits_user_amba_prot_secure(fixer_auto_in_1_a_bits_user_amba_prot_secure),
    .auto_in_1_a_bits_user_amba_prot_fetch(fixer_auto_in_1_a_bits_user_amba_prot_fetch),
    .auto_in_1_a_bits_mask(fixer_auto_in_1_a_bits_mask),
    .auto_in_1_a_bits_data(fixer_auto_in_1_a_bits_data),
    .auto_in_1_d_ready(fixer_auto_in_1_d_ready),
    .auto_in_1_d_valid(fixer_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(fixer_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_size(fixer_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_source(fixer_auto_in_1_d_bits_source),
    .auto_in_1_d_bits_denied(fixer_auto_in_1_d_bits_denied),
    .auto_in_1_d_bits_data(fixer_auto_in_1_d_bits_data),
    .auto_in_1_d_bits_corrupt(fixer_auto_in_1_d_bits_corrupt),
    .auto_in_0_a_ready(fixer_auto_in_0_a_ready),
    .auto_in_0_a_valid(fixer_auto_in_0_a_valid),
    .auto_in_0_a_bits_opcode(fixer_auto_in_0_a_bits_opcode),
    .auto_in_0_a_bits_param(fixer_auto_in_0_a_bits_param),
    .auto_in_0_a_bits_size(fixer_auto_in_0_a_bits_size),
    .auto_in_0_a_bits_source(fixer_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(fixer_auto_in_0_a_bits_address),
    .auto_in_0_a_bits_user_amba_prot_bufferable(fixer_auto_in_0_a_bits_user_amba_prot_bufferable),
    .auto_in_0_a_bits_user_amba_prot_modifiable(fixer_auto_in_0_a_bits_user_amba_prot_modifiable),
    .auto_in_0_a_bits_user_amba_prot_readalloc(fixer_auto_in_0_a_bits_user_amba_prot_readalloc),
    .auto_in_0_a_bits_user_amba_prot_writealloc(fixer_auto_in_0_a_bits_user_amba_prot_writealloc),
    .auto_in_0_a_bits_user_amba_prot_privileged(fixer_auto_in_0_a_bits_user_amba_prot_privileged),
    .auto_in_0_a_bits_user_amba_prot_secure(fixer_auto_in_0_a_bits_user_amba_prot_secure),
    .auto_in_0_a_bits_user_amba_prot_fetch(fixer_auto_in_0_a_bits_user_amba_prot_fetch),
    .auto_in_0_a_bits_mask(fixer_auto_in_0_a_bits_mask),
    .auto_in_0_a_bits_data(fixer_auto_in_0_a_bits_data),
    .auto_in_0_d_ready(fixer_auto_in_0_d_ready),
    .auto_in_0_d_valid(fixer_auto_in_0_d_valid),
    .auto_in_0_d_bits_opcode(fixer_auto_in_0_d_bits_opcode),
    .auto_in_0_d_bits_size(fixer_auto_in_0_d_bits_size),
    .auto_in_0_d_bits_source(fixer_auto_in_0_d_bits_source),
    .auto_in_0_d_bits_denied(fixer_auto_in_0_d_bits_denied),
    .auto_in_0_d_bits_data(fixer_auto_in_0_d_bits_data),
    .auto_in_0_d_bits_corrupt(fixer_auto_in_0_d_bits_corrupt),
    .auto_out_1_a_ready(fixer_auto_out_1_a_ready),
    .auto_out_1_a_valid(fixer_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(fixer_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_param(fixer_auto_out_1_a_bits_param),
    .auto_out_1_a_bits_size(fixer_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(fixer_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(fixer_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_user_amba_prot_bufferable(fixer_auto_out_1_a_bits_user_amba_prot_bufferable),
    .auto_out_1_a_bits_user_amba_prot_modifiable(fixer_auto_out_1_a_bits_user_amba_prot_modifiable),
    .auto_out_1_a_bits_user_amba_prot_readalloc(fixer_auto_out_1_a_bits_user_amba_prot_readalloc),
    .auto_out_1_a_bits_user_amba_prot_writealloc(fixer_auto_out_1_a_bits_user_amba_prot_writealloc),
    .auto_out_1_a_bits_user_amba_prot_privileged(fixer_auto_out_1_a_bits_user_amba_prot_privileged),
    .auto_out_1_a_bits_user_amba_prot_secure(fixer_auto_out_1_a_bits_user_amba_prot_secure),
    .auto_out_1_a_bits_user_amba_prot_fetch(fixer_auto_out_1_a_bits_user_amba_prot_fetch),
    .auto_out_1_a_bits_mask(fixer_auto_out_1_a_bits_mask),
    .auto_out_1_a_bits_data(fixer_auto_out_1_a_bits_data),
    .auto_out_1_d_ready(fixer_auto_out_1_d_ready),
    .auto_out_1_d_valid(fixer_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(fixer_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_size(fixer_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(fixer_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_denied(fixer_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_data(fixer_auto_out_1_d_bits_data),
    .auto_out_1_d_bits_corrupt(fixer_auto_out_1_d_bits_corrupt),
    .auto_out_0_a_ready(fixer_auto_out_0_a_ready),
    .auto_out_0_a_valid(fixer_auto_out_0_a_valid),
    .auto_out_0_a_bits_opcode(fixer_auto_out_0_a_bits_opcode),
    .auto_out_0_a_bits_param(fixer_auto_out_0_a_bits_param),
    .auto_out_0_a_bits_size(fixer_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(fixer_auto_out_0_a_bits_source),
    .auto_out_0_a_bits_address(fixer_auto_out_0_a_bits_address),
    .auto_out_0_a_bits_user_amba_prot_bufferable(fixer_auto_out_0_a_bits_user_amba_prot_bufferable),
    .auto_out_0_a_bits_user_amba_prot_modifiable(fixer_auto_out_0_a_bits_user_amba_prot_modifiable),
    .auto_out_0_a_bits_user_amba_prot_readalloc(fixer_auto_out_0_a_bits_user_amba_prot_readalloc),
    .auto_out_0_a_bits_user_amba_prot_writealloc(fixer_auto_out_0_a_bits_user_amba_prot_writealloc),
    .auto_out_0_a_bits_user_amba_prot_privileged(fixer_auto_out_0_a_bits_user_amba_prot_privileged),
    .auto_out_0_a_bits_user_amba_prot_secure(fixer_auto_out_0_a_bits_user_amba_prot_secure),
    .auto_out_0_a_bits_user_amba_prot_fetch(fixer_auto_out_0_a_bits_user_amba_prot_fetch),
    .auto_out_0_a_bits_mask(fixer_auto_out_0_a_bits_mask),
    .auto_out_0_a_bits_data(fixer_auto_out_0_a_bits_data),
    .auto_out_0_d_ready(fixer_auto_out_0_d_ready),
    .auto_out_0_d_valid(fixer_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(fixer_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_size(fixer_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(fixer_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_denied(fixer_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_data(fixer_auto_out_0_d_bits_data),
    .auto_out_0_d_bits_corrupt(fixer_auto_out_0_d_bits_corrupt),
    .io_covSum(fixer_io_covSum)
  );
  assign subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_clock =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_reset =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_clock =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_reset =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_clock =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_reset =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_clock =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_reset =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_clock =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_reset =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_clock =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_reset =
    subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_clock = clockGroup_auto_in_member_subsystem_sbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_reset = clockGroup_auto_in_member_subsystem_sbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_ready =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_valid =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_opcode =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_size =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_source =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_denied =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_data =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_corrupt =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_valid =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_param =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_size =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_source =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_address =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_mask =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_data =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_ready =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_ready =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_ready; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_valid =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_valid; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_opcode =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_size =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_source =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_denied =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_denied; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_data =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_corrupt =
    coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_valid =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_param =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_size =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_source =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_address =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_mask =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_data =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_ready =
    coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_valid =
    coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_valid; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_opcode =
    coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_param =
    coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_param; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_size =
    coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_source =
    coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_address =
    coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_mask =
    coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_a_bits_data =
    coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_in_d_ready =
    coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_ready; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_a_ready =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_valid =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_opcode =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_size =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_source =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_denied =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_data =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_widget_auto_out_d_bits_corrupt =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_ready =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_valid =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_opcode =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_size =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_source =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_denied =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_data =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_corrupt =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_valid =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_opcode =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_param =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_size =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_source =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_address =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_bufferable =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_modifiable =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_readalloc =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_writealloc =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_privileged =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_secure =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_fetch =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_mask =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_data =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_ready =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_valid =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_valid; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_opcode =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_param =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_param; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_size =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_source =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_address =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_bufferable =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_modifiable =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_readalloc =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_writealloc =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_privileged =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_secure =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_fetch =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_mask =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_data =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_ready =
    coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_ready; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_ready =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_valid =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_opcode =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_size =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_source =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_denied =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_data =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_corrupt =
    coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_valid =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_opcode =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_param =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_size =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_source =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_address =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_bufferable =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_modifiable =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_readalloc =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_writealloc =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_privileged =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_secure =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_user_amba_prot_fetch =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_mask =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_a_bits_data =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_in_d_ready =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_a_ready =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_valid =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_opcode =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_size =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_source =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_denied =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_denied; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_data =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_widget_auto_out_d_bits_corrupt =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_ready =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_d_valid =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_opcode =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_size =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_source =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_denied =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_data =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_corrupt =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_valid =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_size =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_source =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_address =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_bufferable =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_modifiable =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_readalloc =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_writealloc =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_privileged =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_secure =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_fetch =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_mask =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_data =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_d_ready =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_ready =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_a_ready; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_d_valid =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_d_valid; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_opcode =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_size =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_source =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_denied =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_denied; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_data =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_corrupt =
    coupler_to_bus_named_subsystem_l2_widget_auto_in_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_valid =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_size =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_source =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_address =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_bufferable =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_modifiable =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_readalloc =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_writealloc =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_privileged =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_secure =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_fetch =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_mask =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_data =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_ready =
    coupler_to_bus_named_subsystem_l2_widget_auto_out_d_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_valid =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_valid; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_opcode =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_size =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_source =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_address =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_bufferable =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_modifiable =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_readalloc =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_writealloc =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_privileged =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_secure =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_secure; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_user_amba_prot_fetch =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_mask =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_a_bits_data =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_in_d_ready =
    coupler_to_bus_named_subsystem_l2_auto_widget_in_d_ready; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_a_ready =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_d_valid =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_opcode =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_size =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_source =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_denied =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_denied; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_data =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_widget_auto_out_d_bits_corrupt =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_ready = coupler_from_cva6_tile_auto_tl_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_valid = coupler_from_cva6_tile_auto_tl_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_opcode =
    coupler_from_cva6_tile_auto_tl_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_size =
    coupler_from_cva6_tile_auto_tl_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_source =
    coupler_from_cva6_tile_auto_tl_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_denied =
    coupler_from_cva6_tile_auto_tl_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_data =
    coupler_from_cva6_tile_auto_tl_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_corrupt =
    coupler_from_cva6_tile_auto_tl_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_out_a_valid = coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_opcode =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_param =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_size =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_source =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_address =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_bufferable =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_modifiable =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_readalloc =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_writealloc =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_privileged =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_secure =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_fetch =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_mask =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_bits_data =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_d_ready = coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_ready =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_ready; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_valid =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_valid; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_opcode =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_size =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_source =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_denied =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_denied; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_data =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_corrupt =
    coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_bufferable =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_modifiable =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_readalloc =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_writealloc =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_privileged =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_secure =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_fetch =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_ready; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_valid; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_denied; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt =
    coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_param; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_fixedClockNode_out_1_clock = fixedClockNode_auto_out_2_clock; // @[LazyModule.scala 311:12]
  assign auto_fixedClockNode_out_1_reset = fixedClockNode_auto_out_2_reset; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock =
    subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_clock; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset =
    subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_reset; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock =
    subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_clock; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset =
    subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_reset; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock =
    subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_clock; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset =
    subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_reset; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock =
    subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_clock; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset =
    subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_reset; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock =
    subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_clock; // @[LazyModule.scala 311:12]
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset =
    subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_reset; // @[LazyModule.scala 311:12]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock; // @[LazyModule.scala 309:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset; // @[LazyModule.scala 309:16]
  assign clockGroup_auto_in_member_subsystem_sbus_0_clock =
    subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_clock; // @[LazyModule.scala 298:16]
  assign clockGroup_auto_in_member_subsystem_sbus_0_reset =
    subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_reset; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign system_bus_xbar_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_valid = fixer_auto_out_1_a_valid; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_opcode = fixer_auto_out_1_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_param = fixer_auto_out_1_a_bits_param; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_size = fixer_auto_out_1_a_bits_size; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_source = fixer_auto_out_1_a_bits_source; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_address = fixer_auto_out_1_a_bits_address; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_user_amba_prot_bufferable = fixer_auto_out_1_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_user_amba_prot_modifiable = fixer_auto_out_1_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_user_amba_prot_readalloc = fixer_auto_out_1_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_user_amba_prot_writealloc = fixer_auto_out_1_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_user_amba_prot_privileged = fixer_auto_out_1_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_user_amba_prot_secure = fixer_auto_out_1_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_user_amba_prot_fetch = fixer_auto_out_1_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_mask = fixer_auto_out_1_a_bits_mask; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_a_bits_data = fixer_auto_out_1_a_bits_data; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_1_d_ready = fixer_auto_out_1_d_ready; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_valid = fixer_auto_out_0_a_valid; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_opcode = fixer_auto_out_0_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_param = fixer_auto_out_0_a_bits_param; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_size = fixer_auto_out_0_a_bits_size; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_source = fixer_auto_out_0_a_bits_source; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_address = fixer_auto_out_0_a_bits_address; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_user_amba_prot_bufferable = fixer_auto_out_0_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_user_amba_prot_modifiable = fixer_auto_out_0_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_user_amba_prot_readalloc = fixer_auto_out_0_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_user_amba_prot_writealloc = fixer_auto_out_0_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_user_amba_prot_privileged = fixer_auto_out_0_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_user_amba_prot_secure = fixer_auto_out_0_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_user_amba_prot_fetch = fixer_auto_out_0_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_mask = fixer_auto_out_0_a_bits_mask; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_a_bits_data = fixer_auto_out_0_a_bits_data; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_in_0_d_ready = fixer_auto_out_0_d_ready; // @[LazyModule.scala 296:16]
  assign system_bus_xbar_auto_out_1_a_ready = coupler_to_bus_named_subsystem_l2_auto_widget_in_a_ready; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_1_d_valid = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_valid; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_1_d_bits_opcode = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_1_d_bits_size = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_1_d_bits_source = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_1_d_bits_denied = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_1_d_bits_data = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_1_d_bits_corrupt = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_0_a_ready = coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_ready; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_0_d_valid = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_valid; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_0_d_bits_opcode = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_0_d_bits_size = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_0_d_bits_source = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_0_d_bits_denied = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_0_d_bits_data = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign system_bus_xbar_auto_out_0_d_bits_corrupt = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign fixer_auto_in_1_a_valid = coupler_from_cva6_tile_auto_tl_out_a_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_opcode = coupler_from_cva6_tile_auto_tl_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_param = coupler_from_cva6_tile_auto_tl_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_size = coupler_from_cva6_tile_auto_tl_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_source = coupler_from_cva6_tile_auto_tl_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_address = coupler_from_cva6_tile_auto_tl_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_user_amba_prot_bufferable =
    coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_user_amba_prot_modifiable =
    coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_user_amba_prot_readalloc =
    coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_user_amba_prot_writealloc =
    coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_user_amba_prot_privileged =
    coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_user_amba_prot_secure = coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_user_amba_prot_fetch = coupler_from_cva6_tile_auto_tl_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_mask = coupler_from_cva6_tile_auto_tl_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_a_bits_data = coupler_from_cva6_tile_auto_tl_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_1_d_ready = coupler_from_cva6_tile_auto_tl_out_d_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_valid = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_opcode = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_param = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_size = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_source = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_address = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_user_amba_prot_bufferable =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_user_amba_prot_modifiable =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_user_amba_prot_readalloc =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_user_amba_prot_writealloc =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_user_amba_prot_privileged =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_user_amba_prot_secure =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_user_amba_prot_fetch =
    coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_mask = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_a_bits_data = coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_0_d_ready = coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_1_a_ready = system_bus_xbar_auto_in_1_a_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_1_d_valid = system_bus_xbar_auto_in_1_d_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_1_d_bits_opcode = system_bus_xbar_auto_in_1_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_1_d_bits_size = system_bus_xbar_auto_in_1_d_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_1_d_bits_source = system_bus_xbar_auto_in_1_d_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_1_d_bits_denied = system_bus_xbar_auto_in_1_d_bits_denied; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_1_d_bits_data = system_bus_xbar_auto_in_1_d_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_1_d_bits_corrupt = system_bus_xbar_auto_in_1_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_0_a_ready = system_bus_xbar_auto_in_0_a_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_0_d_valid = system_bus_xbar_auto_in_0_d_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_0_d_bits_opcode = system_bus_xbar_auto_in_0_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_0_d_bits_size = system_bus_xbar_auto_in_0_d_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_0_d_bits_source = system_bus_xbar_auto_in_0_d_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_0_d_bits_denied = system_bus_xbar_auto_in_0_d_bits_denied; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_0_d_bits_data = system_bus_xbar_auto_in_0_d_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_0_d_bits_corrupt = system_bus_xbar_auto_in_0_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_valid = system_bus_xbar_auto_out_0_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_opcode = system_bus_xbar_auto_out_0_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_param = system_bus_xbar_auto_out_0_a_bits_param; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_size = system_bus_xbar_auto_out_0_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_source = system_bus_xbar_auto_out_0_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_address = system_bus_xbar_auto_out_0_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_mask = system_bus_xbar_auto_out_0_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_data = system_bus_xbar_auto_out_0_a_bits_data; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_ready = system_bus_xbar_auto_out_0_d_ready; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_ready =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_valid =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_opcode =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_size =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_source =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_denied =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_data =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_corrupt =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_a_ready = fixer_auto_in_0_a_ready; // @[LazyModule.scala 296:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_valid = fixer_auto_in_0_d_valid; // @[LazyModule.scala 296:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_opcode = fixer_auto_in_0_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_size = fixer_auto_in_0_d_bits_size; // @[LazyModule.scala 296:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_source = fixer_auto_in_0_d_bits_source; // @[LazyModule.scala 296:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_denied = fixer_auto_in_0_d_bits_denied; // @[LazyModule.scala 296:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_data = fixer_auto_in_0_d_bits_data; // @[LazyModule.scala 296:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_widget_out_d_bits_corrupt = fixer_auto_in_0_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_valid =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_opcode =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_param =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_size =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_source =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_address =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_bufferable =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_modifiable =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_readalloc =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_writealloc =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_privileged =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_secure =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_secure; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_user_amba_prot_fetch =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_mask =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_a_bits_data =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_from_bus_named_subsystem_fbus_auto_bus_xing_in_d_ready =
    auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_valid = system_bus_xbar_auto_out_1_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_opcode = system_bus_xbar_auto_out_1_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_size = system_bus_xbar_auto_out_1_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_source = system_bus_xbar_auto_out_1_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_address = system_bus_xbar_auto_out_1_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_bufferable =
    system_bus_xbar_auto_out_1_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_modifiable =
    system_bus_xbar_auto_out_1_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_readalloc =
    system_bus_xbar_auto_out_1_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_writealloc =
    system_bus_xbar_auto_out_1_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_privileged =
    system_bus_xbar_auto_out_1_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_secure =
    system_bus_xbar_auto_out_1_a_bits_user_amba_prot_secure; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_user_amba_prot_fetch =
    system_bus_xbar_auto_out_1_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_mask = system_bus_xbar_auto_out_1_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_data = system_bus_xbar_auto_out_1_a_bits_data; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_d_ready = system_bus_xbar_auto_out_1_d_ready; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_ready =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_valid =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_opcode =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_size =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_source =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_denied =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_data =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_corrupt =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_valid =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_valid; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_opcode =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_param =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_param; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_size =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_source =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_address =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_bufferable =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_modifiable =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_readalloc =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_writealloc =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_privileged =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_secure =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_secure; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_user_amba_prot_fetch =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_mask =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_a_bits_data =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_master_clock_xing_in_d_ready =
    auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_ready; // @[LazyModule.scala 309:16]
  assign coupler_from_cva6_tile_auto_tl_out_a_ready = fixer_auto_in_1_a_ready; // @[LazyModule.scala 296:16]
  assign coupler_from_cva6_tile_auto_tl_out_d_valid = fixer_auto_in_1_d_valid; // @[LazyModule.scala 296:16]
  assign coupler_from_cva6_tile_auto_tl_out_d_bits_opcode = fixer_auto_in_1_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign coupler_from_cva6_tile_auto_tl_out_d_bits_size = fixer_auto_in_1_d_bits_size; // @[LazyModule.scala 296:16]
  assign coupler_from_cva6_tile_auto_tl_out_d_bits_source = fixer_auto_in_1_d_bits_source; // @[LazyModule.scala 296:16]
  assign coupler_from_cva6_tile_auto_tl_out_d_bits_denied = fixer_auto_in_1_d_bits_denied; // @[LazyModule.scala 296:16]
  assign coupler_from_cva6_tile_auto_tl_out_d_bits_data = fixer_auto_in_1_d_bits_data; // @[LazyModule.scala 296:16]
  assign coupler_from_cva6_tile_auto_tl_out_d_bits_corrupt = fixer_auto_in_1_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign SystemBus_covSum = 30'h0;
  assign fixedClockNode_sum = SystemBus_covSum + fixedClockNode_io_covSum;
  assign system_bus_xbar_sum = fixedClockNode_sum + system_bus_xbar_io_covSum;
  assign fixer_sum = system_bus_xbar_sum + fixer_io_covSum;
  assign io_covSum = fixer_sum;
  assign system_bus_xbar_metaReset = metaReset;
endmodule
module FixedClockBroadcast_1(
  input         auto_in_clock,
  input         auto_in_reset,
  output        auto_out_1_clock,
  output        auto_out_1_reset,
  output        auto_out_0_clock,
  output        auto_out_0_reset,
  output [29:0] io_covSum
);
  wire [29:0] FixedClockBroadcast_1_covSum;
  assign auto_out_1_clock = auto_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_reset = auto_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_clock = auto_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_reset = auto_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign FixedClockBroadcast_1_covSum = 30'h0;
  assign io_covSum = FixedClockBroadcast_1_covSum;
endmodule
module TLFIFOFixer_1(
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [30:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [30:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [2:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input  [63:0] auto_out_d_bits_data,
  output [29:0] io_covSum
);
  wire [29:0] TLFIFOFixer_1_covSum;
  assign auto_in_a_ready = auto_out_a_ready; // @[FIFOFixer.scala 88:33]
  assign auto_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[FIFOFixer.scala 87:33]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLFIFOFixer_1_covSum = 30'h0;
  assign io_covSum = TLFIFOFixer_1_covSum;
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [30:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [30:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_param_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [6:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg [30:0] ram_address [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [30:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [30:0] ram_address_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_en = 1'h1;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_covSum = 30'h0;
  assign io_covSum = Queue_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= value_1 + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  value_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input         io_enq_bits_denied,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output        io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [6:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_denied [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_1_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_1_covSum = 30'h0;
  assign io_covSum = Queue_1_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= value_1 + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_5[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  value_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [30:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [2:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [30:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [2:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum
);
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_param; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire [30:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 361:21]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [30:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 361:21]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [29:0] bundleOut_0_a_q_io_covSum; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire [29:0] bundleIn_0_d_q_io_covSum; // @[Decoupled.scala 361:21]
  wire [29:0] TLBuffer_covSum;
  wire [29:0] bundleOut_0_a_q_sum;
  wire [29:0] bundleIn_0_d_q_sum;
  Queue bundleOut_0_a_q ( // @[Decoupled.scala 361:21]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_covSum(bundleOut_0_a_q_io_covSum)
  );
  Queue_1 bundleIn_0_d_q ( // @[Decoupled.scala 361:21]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt),
    .io_covSum(bundleIn_0_d_q_io_covSum)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 Decoupled.scala 365:17]
  assign bundleOut_0_a_q_clock = clock;
  assign bundleOut_0_a_q_reset = reset;
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_clock = clock;
  assign bundleIn_0_d_q_reset = reset;
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBuffer_covSum = 30'h0;
  assign bundleOut_0_a_q_sum = TLBuffer_covSum + bundleOut_0_a_q_io_covSum;
  assign bundleIn_0_d_q_sum = bundleOut_0_a_q_sum + bundleIn_0_d_q_io_covSum;
  assign io_covSum = bundleIn_0_d_q_sum;
endmodule
module TLAtomicAutomata(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [30:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [2:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [30:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [2:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] cam_s_0_state; // @[AtomicAutomata.scala 76:28]
  reg [2:0] cam_a_0_bits_opcode; // @[AtomicAutomata.scala 77:24]
  reg [2:0] cam_a_0_bits_param; // @[AtomicAutomata.scala 77:24]
  reg [2:0] cam_a_0_bits_size; // @[AtomicAutomata.scala 77:24]
  reg [6:0] cam_a_0_bits_source; // @[AtomicAutomata.scala 77:24]
  reg [30:0] cam_a_0_bits_address; // @[AtomicAutomata.scala 77:24]
  reg [7:0] cam_a_0_bits_mask; // @[AtomicAutomata.scala 77:24]
  reg [63:0] cam_a_0_bits_data; // @[AtomicAutomata.scala 77:24]
  reg [3:0] cam_a_0_lut; // @[AtomicAutomata.scala 77:24]
  reg [63:0] cam_d_0_data; // @[AtomicAutomata.scala 78:24]
  reg  cam_d_0_denied; // @[AtomicAutomata.scala 78:24]
  reg  cam_d_0_corrupt; // @[AtomicAutomata.scala 78:24]
  wire  cam_free_0 = cam_s_0_state == 2'h0; // @[AtomicAutomata.scala 80:44]
  wire  cam_amo_0 = cam_s_0_state == 2'h2; // @[AtomicAutomata.scala 81:44]
  wire  cam_abusy_0 = cam_s_0_state == 2'h3 | cam_amo_0; // @[AtomicAutomata.scala 82:57]
  wire  cam_dmatch_0 = cam_s_0_state != 2'h0; // @[AtomicAutomata.scala 83:49]
  wire  a_isLogical = auto_in_a_bits_opcode == 3'h3; // @[AtomicAutomata.scala 90:47]
  wire  a_isArithmetic = auto_in_a_bits_opcode == 3'h2; // @[AtomicAutomata.scala 91:47]
  wire  _a_isSupported_T = a_isArithmetic ? 1'h0 : 1'h1; // @[AtomicAutomata.scala 92:63]
  wire  a_isSupported = a_isLogical ? 1'h0 : _a_isSupported_T; // @[AtomicAutomata.scala 92:32]
  wire [1:0] indexes_0 = {cam_a_0_bits_data[0],cam_d_0_data[0]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_1 = {cam_a_0_bits_data[1],cam_d_0_data[1]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_2 = {cam_a_0_bits_data[2],cam_d_0_data[2]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_3 = {cam_a_0_bits_data[3],cam_d_0_data[3]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_4 = {cam_a_0_bits_data[4],cam_d_0_data[4]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_5 = {cam_a_0_bits_data[5],cam_d_0_data[5]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_6 = {cam_a_0_bits_data[6],cam_d_0_data[6]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_7 = {cam_a_0_bits_data[7],cam_d_0_data[7]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_8 = {cam_a_0_bits_data[8],cam_d_0_data[8]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_9 = {cam_a_0_bits_data[9],cam_d_0_data[9]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_10 = {cam_a_0_bits_data[10],cam_d_0_data[10]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_11 = {cam_a_0_bits_data[11],cam_d_0_data[11]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_12 = {cam_a_0_bits_data[12],cam_d_0_data[12]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_13 = {cam_a_0_bits_data[13],cam_d_0_data[13]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_14 = {cam_a_0_bits_data[14],cam_d_0_data[14]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_15 = {cam_a_0_bits_data[15],cam_d_0_data[15]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_16 = {cam_a_0_bits_data[16],cam_d_0_data[16]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_17 = {cam_a_0_bits_data[17],cam_d_0_data[17]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_18 = {cam_a_0_bits_data[18],cam_d_0_data[18]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_19 = {cam_a_0_bits_data[19],cam_d_0_data[19]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_20 = {cam_a_0_bits_data[20],cam_d_0_data[20]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_21 = {cam_a_0_bits_data[21],cam_d_0_data[21]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_22 = {cam_a_0_bits_data[22],cam_d_0_data[22]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_23 = {cam_a_0_bits_data[23],cam_d_0_data[23]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_24 = {cam_a_0_bits_data[24],cam_d_0_data[24]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_25 = {cam_a_0_bits_data[25],cam_d_0_data[25]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_26 = {cam_a_0_bits_data[26],cam_d_0_data[26]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_27 = {cam_a_0_bits_data[27],cam_d_0_data[27]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_28 = {cam_a_0_bits_data[28],cam_d_0_data[28]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_29 = {cam_a_0_bits_data[29],cam_d_0_data[29]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_30 = {cam_a_0_bits_data[30],cam_d_0_data[30]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_31 = {cam_a_0_bits_data[31],cam_d_0_data[31]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_32 = {cam_a_0_bits_data[32],cam_d_0_data[32]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_33 = {cam_a_0_bits_data[33],cam_d_0_data[33]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_34 = {cam_a_0_bits_data[34],cam_d_0_data[34]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_35 = {cam_a_0_bits_data[35],cam_d_0_data[35]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_36 = {cam_a_0_bits_data[36],cam_d_0_data[36]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_37 = {cam_a_0_bits_data[37],cam_d_0_data[37]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_38 = {cam_a_0_bits_data[38],cam_d_0_data[38]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_39 = {cam_a_0_bits_data[39],cam_d_0_data[39]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_40 = {cam_a_0_bits_data[40],cam_d_0_data[40]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_41 = {cam_a_0_bits_data[41],cam_d_0_data[41]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_42 = {cam_a_0_bits_data[42],cam_d_0_data[42]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_43 = {cam_a_0_bits_data[43],cam_d_0_data[43]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_44 = {cam_a_0_bits_data[44],cam_d_0_data[44]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_45 = {cam_a_0_bits_data[45],cam_d_0_data[45]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_46 = {cam_a_0_bits_data[46],cam_d_0_data[46]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_47 = {cam_a_0_bits_data[47],cam_d_0_data[47]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_48 = {cam_a_0_bits_data[48],cam_d_0_data[48]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_49 = {cam_a_0_bits_data[49],cam_d_0_data[49]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_50 = {cam_a_0_bits_data[50],cam_d_0_data[50]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_51 = {cam_a_0_bits_data[51],cam_d_0_data[51]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_52 = {cam_a_0_bits_data[52],cam_d_0_data[52]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_53 = {cam_a_0_bits_data[53],cam_d_0_data[53]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_54 = {cam_a_0_bits_data[54],cam_d_0_data[54]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_55 = {cam_a_0_bits_data[55],cam_d_0_data[55]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_56 = {cam_a_0_bits_data[56],cam_d_0_data[56]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_57 = {cam_a_0_bits_data[57],cam_d_0_data[57]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_58 = {cam_a_0_bits_data[58],cam_d_0_data[58]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_59 = {cam_a_0_bits_data[59],cam_d_0_data[59]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_60 = {cam_a_0_bits_data[60],cam_d_0_data[60]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_61 = {cam_a_0_bits_data[61],cam_d_0_data[61]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_62 = {cam_a_0_bits_data[62],cam_d_0_data[62]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_63 = {cam_a_0_bits_data[63],cam_d_0_data[63]}; // @[Cat.scala 31:58]
  wire [3:0] _logic_out_T = cam_a_0_lut >> indexes_0; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_2 = cam_a_0_lut >> indexes_1; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_4 = cam_a_0_lut >> indexes_2; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_6 = cam_a_0_lut >> indexes_3; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_8 = cam_a_0_lut >> indexes_4; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_10 = cam_a_0_lut >> indexes_5; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_12 = cam_a_0_lut >> indexes_6; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_14 = cam_a_0_lut >> indexes_7; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_16 = cam_a_0_lut >> indexes_8; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_18 = cam_a_0_lut >> indexes_9; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_20 = cam_a_0_lut >> indexes_10; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_22 = cam_a_0_lut >> indexes_11; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_24 = cam_a_0_lut >> indexes_12; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_26 = cam_a_0_lut >> indexes_13; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_28 = cam_a_0_lut >> indexes_14; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_30 = cam_a_0_lut >> indexes_15; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_32 = cam_a_0_lut >> indexes_16; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_34 = cam_a_0_lut >> indexes_17; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_36 = cam_a_0_lut >> indexes_18; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_38 = cam_a_0_lut >> indexes_19; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_40 = cam_a_0_lut >> indexes_20; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_42 = cam_a_0_lut >> indexes_21; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_44 = cam_a_0_lut >> indexes_22; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_46 = cam_a_0_lut >> indexes_23; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_48 = cam_a_0_lut >> indexes_24; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_50 = cam_a_0_lut >> indexes_25; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_52 = cam_a_0_lut >> indexes_26; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_54 = cam_a_0_lut >> indexes_27; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_56 = cam_a_0_lut >> indexes_28; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_58 = cam_a_0_lut >> indexes_29; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_60 = cam_a_0_lut >> indexes_30; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_62 = cam_a_0_lut >> indexes_31; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_64 = cam_a_0_lut >> indexes_32; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_66 = cam_a_0_lut >> indexes_33; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_68 = cam_a_0_lut >> indexes_34; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_70 = cam_a_0_lut >> indexes_35; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_72 = cam_a_0_lut >> indexes_36; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_74 = cam_a_0_lut >> indexes_37; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_76 = cam_a_0_lut >> indexes_38; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_78 = cam_a_0_lut >> indexes_39; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_80 = cam_a_0_lut >> indexes_40; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_82 = cam_a_0_lut >> indexes_41; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_84 = cam_a_0_lut >> indexes_42; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_86 = cam_a_0_lut >> indexes_43; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_88 = cam_a_0_lut >> indexes_44; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_90 = cam_a_0_lut >> indexes_45; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_92 = cam_a_0_lut >> indexes_46; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_94 = cam_a_0_lut >> indexes_47; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_96 = cam_a_0_lut >> indexes_48; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_98 = cam_a_0_lut >> indexes_49; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_100 = cam_a_0_lut >> indexes_50; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_102 = cam_a_0_lut >> indexes_51; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_104 = cam_a_0_lut >> indexes_52; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_106 = cam_a_0_lut >> indexes_53; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_108 = cam_a_0_lut >> indexes_54; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_110 = cam_a_0_lut >> indexes_55; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_112 = cam_a_0_lut >> indexes_56; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_114 = cam_a_0_lut >> indexes_57; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_116 = cam_a_0_lut >> indexes_58; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_118 = cam_a_0_lut >> indexes_59; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_120 = cam_a_0_lut >> indexes_60; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_122 = cam_a_0_lut >> indexes_61; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_124 = cam_a_0_lut >> indexes_62; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_126 = cam_a_0_lut >> indexes_63; // @[AtomicAutomata.scala 114:57]
  wire [7:0] logic_out_lo_lo_lo = {_logic_out_T_14[0],_logic_out_T_12[0],_logic_out_T_10[0],_logic_out_T_8[0],
    _logic_out_T_6[0],_logic_out_T_4[0],_logic_out_T_2[0],_logic_out_T[0]}; // @[Cat.scala 31:58]
  wire [15:0] logic_out_lo_lo = {_logic_out_T_30[0],_logic_out_T_28[0],_logic_out_T_26[0],_logic_out_T_24[0],
    _logic_out_T_22[0],_logic_out_T_20[0],_logic_out_T_18[0],_logic_out_T_16[0],logic_out_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] logic_out_lo_hi_lo = {_logic_out_T_46[0],_logic_out_T_44[0],_logic_out_T_42[0],_logic_out_T_40[0],
    _logic_out_T_38[0],_logic_out_T_36[0],_logic_out_T_34[0],_logic_out_T_32[0]}; // @[Cat.scala 31:58]
  wire [31:0] logic_out_lo = {_logic_out_T_62[0],_logic_out_T_60[0],_logic_out_T_58[0],_logic_out_T_56[0],
    _logic_out_T_54[0],_logic_out_T_52[0],_logic_out_T_50[0],_logic_out_T_48[0],logic_out_lo_hi_lo,logic_out_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] logic_out_hi_lo_lo = {_logic_out_T_78[0],_logic_out_T_76[0],_logic_out_T_74[0],_logic_out_T_72[0],
    _logic_out_T_70[0],_logic_out_T_68[0],_logic_out_T_66[0],_logic_out_T_64[0]}; // @[Cat.scala 31:58]
  wire [15:0] logic_out_hi_lo = {_logic_out_T_94[0],_logic_out_T_92[0],_logic_out_T_90[0],_logic_out_T_88[0],
    _logic_out_T_86[0],_logic_out_T_84[0],_logic_out_T_82[0],_logic_out_T_80[0],logic_out_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] logic_out_hi_hi_lo = {_logic_out_T_110[0],_logic_out_T_108[0],_logic_out_T_106[0],_logic_out_T_104[0],
    _logic_out_T_102[0],_logic_out_T_100[0],_logic_out_T_98[0],_logic_out_T_96[0]}; // @[Cat.scala 31:58]
  wire [31:0] logic_out_hi = {_logic_out_T_126[0],_logic_out_T_124[0],_logic_out_T_122[0],_logic_out_T_120[0],
    _logic_out_T_118[0],_logic_out_T_116[0],_logic_out_T_114[0],_logic_out_T_112[0],logic_out_hi_hi_lo,logic_out_hi_lo}; // @[Cat.scala 31:58]
  wire [63:0] logic_out = {logic_out_hi,logic_out_lo}; // @[Cat.scala 31:58]
  wire  unsigned_ = cam_a_0_bits_param[1]; // @[AtomicAutomata.scala 117:42]
  wire  take_max = cam_a_0_bits_param[0]; // @[AtomicAutomata.scala 118:42]
  wire  adder = cam_a_0_bits_param[2]; // @[AtomicAutomata.scala 119:39]
  wire [7:0] _signSel_T = ~cam_a_0_bits_mask; // @[AtomicAutomata.scala 121:25]
  wire [7:0] _GEN_10 = {{1'd0}, cam_a_0_bits_mask[7:1]}; // @[AtomicAutomata.scala 121:31]
  wire [7:0] _signSel_T_2 = _signSel_T | _GEN_10; // @[AtomicAutomata.scala 121:31]
  wire [7:0] signSel = ~_signSel_T_2; // @[AtomicAutomata.scala 121:23]
  wire [7:0] signbits_a = {cam_a_0_bits_data[63],cam_a_0_bits_data[55],cam_a_0_bits_data[47],cam_a_0_bits_data[39],
    cam_a_0_bits_data[31],cam_a_0_bits_data[23],cam_a_0_bits_data[15],cam_a_0_bits_data[7]}; // @[Cat.scala 31:58]
  wire [7:0] signbits_d = {cam_d_0_data[63],cam_d_0_data[55],cam_d_0_data[47],cam_d_0_data[39],cam_d_0_data[31],
    cam_d_0_data[23],cam_d_0_data[15],cam_d_0_data[7]}; // @[Cat.scala 31:58]
  wire [7:0] _signbit_a_T = signbits_a & signSel; // @[AtomicAutomata.scala 125:38]
  wire [8:0] _signbit_a_T_1 = {_signbit_a_T, 1'h0}; // @[AtomicAutomata.scala 125:49]
  wire [7:0] signbit_a = _signbit_a_T_1[7:0]; // @[AtomicAutomata.scala 125:54]
  wire [7:0] _signbit_d_T = signbits_d & signSel; // @[AtomicAutomata.scala 126:38]
  wire [8:0] _signbit_d_T_1 = {_signbit_d_T, 1'h0}; // @[AtomicAutomata.scala 126:49]
  wire [7:0] signbit_d = _signbit_d_T_1[7:0]; // @[AtomicAutomata.scala 126:54]
  wire [8:0] _signext_a_T = {signbit_a, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_a_T_2 = signbit_a | _signext_a_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _signext_a_T_3 = {_signext_a_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_a_T_5 = _signext_a_T_2 | _signext_a_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _signext_a_T_6 = {_signext_a_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_a_T_8 = _signext_a_T_5 | _signext_a_T_6[7:0]; // @[package.scala 244:43]
  wire [7:0] _signext_a_T_19 = _signext_a_T_8[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_21 = _signext_a_T_8[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_23 = _signext_a_T_8[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_25 = _signext_a_T_8[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_27 = _signext_a_T_8[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_29 = _signext_a_T_8[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_31 = _signext_a_T_8[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_33 = _signext_a_T_8[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] signext_a = {_signext_a_T_33,_signext_a_T_31,_signext_a_T_29,_signext_a_T_27,_signext_a_T_25,
    _signext_a_T_23,_signext_a_T_21,_signext_a_T_19}; // @[Cat.scala 31:58]
  wire [8:0] _signext_d_T = {signbit_d, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_d_T_2 = signbit_d | _signext_d_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _signext_d_T_3 = {_signext_d_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_d_T_5 = _signext_d_T_2 | _signext_d_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _signext_d_T_6 = {_signext_d_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_d_T_8 = _signext_d_T_5 | _signext_d_T_6[7:0]; // @[package.scala 244:43]
  wire [7:0] _signext_d_T_19 = _signext_d_T_8[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_21 = _signext_d_T_8[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_23 = _signext_d_T_8[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_25 = _signext_d_T_8[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_27 = _signext_d_T_8[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_29 = _signext_d_T_8[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_31 = _signext_d_T_8[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_33 = _signext_d_T_8[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] signext_d = {_signext_d_T_33,_signext_d_T_31,_signext_d_T_29,_signext_d_T_27,_signext_d_T_25,
    _signext_d_T_23,_signext_d_T_21,_signext_d_T_19}; // @[Cat.scala 31:58]
  wire [7:0] _wide_mask_T_9 = cam_a_0_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_11 = cam_a_0_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_13 = cam_a_0_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_15 = cam_a_0_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_17 = cam_a_0_bits_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_19 = cam_a_0_bits_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_21 = cam_a_0_bits_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_23 = cam_a_0_bits_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] wide_mask = {_wide_mask_T_23,_wide_mask_T_21,_wide_mask_T_19,_wide_mask_T_17,_wide_mask_T_15,
    _wide_mask_T_13,_wide_mask_T_11,_wide_mask_T_9}; // @[Cat.scala 31:58]
  wire [63:0] _a_a_ext_T = cam_a_0_bits_data & wide_mask; // @[AtomicAutomata.scala 131:28]
  wire [63:0] a_a_ext = _a_a_ext_T | signext_a; // @[AtomicAutomata.scala 131:41]
  wire [63:0] _a_d_ext_T = cam_d_0_data & wide_mask; // @[AtomicAutomata.scala 132:28]
  wire [63:0] a_d_ext = _a_d_ext_T | signext_d; // @[AtomicAutomata.scala 132:41]
  wire [63:0] _a_d_inv_T = ~a_d_ext; // @[AtomicAutomata.scala 133:43]
  wire [63:0] a_d_inv = adder ? a_d_ext : _a_d_inv_T; // @[AtomicAutomata.scala 133:26]
  wire [63:0] adder_out = a_a_ext + a_d_inv; // @[AtomicAutomata.scala 134:33]
  wire  a_bigger_uneq = unsigned_ == a_a_ext[63]; // @[AtomicAutomata.scala 136:38]
  wire  a_bigger = a_a_ext[63] == a_d_ext[63] ? ~adder_out[63] : a_bigger_uneq; // @[AtomicAutomata.scala 137:27]
  wire  pick_a = take_max == a_bigger; // @[AtomicAutomata.scala 138:31]
  wire [63:0] _arith_out_T = pick_a ? cam_a_0_bits_data : cam_d_0_data; // @[AtomicAutomata.scala 139:50]
  wire [63:0] arith_out = adder ? adder_out : _arith_out_T; // @[AtomicAutomata.scala 139:28]
  wire [63:0] amo_data = cam_a_0_bits_opcode[0] ? logic_out : arith_out; // @[AtomicAutomata.scala 145:14]
  wire  a_allow = ~cam_abusy_0 & (a_isSupported | cam_free_0); // @[AtomicAutomata.scala 149:35]
  reg [2:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 3'h0; // @[Arbiter.scala 88:28]
  wire  source_i_valid = auto_in_a_valid & a_allow; // @[AtomicAutomata.scala 151:38]
  wire [1:0] _readys_T = {source_i_valid,cam_amo_0}; // @[Cat.scala 31:58]
  wire [2:0] _readys_T_1 = {_readys_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0]; // @[package.scala 244:43]
  wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0}; // @[Arbiter.scala 16:78]
  wire [1:0] _readys_T_7 = ~_readys_T_5[1:0]; // @[Arbiter.scala 16:61]
  wire  readys_1 = _readys_T_7[1]; // @[Arbiter.scala 95:86]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 123:31]
  wire  _T = ~a_isSupported; // @[AtomicAutomata.scala 153:15]
  wire [2:0] source_i_bits_opcode = ~a_isSupported ? 3'h4 : auto_in_a_bits_opcode; // @[AtomicAutomata.scala 152:24 153:31 154:32]
  wire [2:0] source_i_bits_param = ~a_isSupported ? 3'h0 : auto_in_a_bits_param; // @[AtomicAutomata.scala 152:24 153:31 155:32]
  wire [1:0] source_c_bits_a_mask_sizeOH_shiftAmount = cam_a_0_bits_size[1:0]; // @[OneHot.scala 63:49]
  wire [3:0] _source_c_bits_a_mask_sizeOH_T_1 = 4'h1 << source_c_bits_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [2:0] source_c_bits_a_mask_sizeOH = _source_c_bits_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _source_c_bits_a_mask_T = cam_a_0_bits_size >= 3'h3; // @[Misc.scala 205:21]
  wire  source_c_bits_a_mask_size = source_c_bits_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  source_c_bits_a_mask_bit = cam_a_0_bits_address[2]; // @[Misc.scala 209:26]
  wire  source_c_bits_a_mask_nbit = ~source_c_bits_a_mask_bit; // @[Misc.scala 210:20]
  wire  source_c_bits_a_mask_acc = _source_c_bits_a_mask_T | source_c_bits_a_mask_size & source_c_bits_a_mask_nbit; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_acc_1 = _source_c_bits_a_mask_T | source_c_bits_a_mask_size & source_c_bits_a_mask_bit; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_size_1 = source_c_bits_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  source_c_bits_a_mask_bit_1 = cam_a_0_bits_address[1]; // @[Misc.scala 209:26]
  wire  source_c_bits_a_mask_nbit_1 = ~source_c_bits_a_mask_bit_1; // @[Misc.scala 210:20]
  wire  source_c_bits_a_mask_eq_2 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_2 = source_c_bits_a_mask_acc | source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_2; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_3 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_3 = source_c_bits_a_mask_acc | source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_3; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_4 = source_c_bits_a_mask_bit & source_c_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_4 = source_c_bits_a_mask_acc_1 | source_c_bits_a_mask_size_1 &
    source_c_bits_a_mask_eq_4; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_5 = source_c_bits_a_mask_bit & source_c_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_5 = source_c_bits_a_mask_acc_1 | source_c_bits_a_mask_size_1 &
    source_c_bits_a_mask_eq_5; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_size_2 = source_c_bits_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  source_c_bits_a_mask_bit_2 = cam_a_0_bits_address[0]; // @[Misc.scala 209:26]
  wire  source_c_bits_a_mask_nbit_2 = ~source_c_bits_a_mask_bit_2; // @[Misc.scala 210:20]
  wire  source_c_bits_a_mask_eq_6 = source_c_bits_a_mask_eq_2 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_6 = source_c_bits_a_mask_acc_2 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_6; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_7 = source_c_bits_a_mask_eq_2 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_7 = source_c_bits_a_mask_acc_2 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_7; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_8 = source_c_bits_a_mask_eq_3 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_8 = source_c_bits_a_mask_acc_3 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_8; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_9 = source_c_bits_a_mask_eq_3 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_9 = source_c_bits_a_mask_acc_3 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_9; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_10 = source_c_bits_a_mask_eq_4 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_10 = source_c_bits_a_mask_acc_4 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_10; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_11 = source_c_bits_a_mask_eq_4 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_11 = source_c_bits_a_mask_acc_4 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_11; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_12 = source_c_bits_a_mask_eq_5 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_12 = source_c_bits_a_mask_acc_5 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_12; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_13 = source_c_bits_a_mask_eq_5 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_13 = source_c_bits_a_mask_acc_5 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] source_c_bits_a_mask = {source_c_bits_a_mask_acc_13,source_c_bits_a_mask_acc_12,source_c_bits_a_mask_acc_11
    ,source_c_bits_a_mask_acc_10,source_c_bits_a_mask_acc_9,source_c_bits_a_mask_acc_8,source_c_bits_a_mask_acc_7,
    source_c_bits_a_mask_acc_6}; // @[Cat.scala 31:58]
  wire [12:0] _decode_T_1 = 13'h3f << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _decode_T_3 = ~_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] decode = _decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 89:24]
  wire  readys_0 = _readys_T_7[0]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_0 = readys_0 & cam_amo_0; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1 = readys_1 & source_i_valid; // @[Arbiter.scala 97:79]
  wire  _T_10 = ~reset; // @[Arbiter.scala 105:13]
  wire  _T_12 = cam_amo_0 | source_i_valid; // @[Arbiter.scala 107:36]
  wire  _T_13 = ~(cam_amo_0 | source_i_valid); // @[Arbiter.scala 107:15]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & cam_amo_0 | state_1 & source_i_valid; // @[Mux.scala 27:73]
  wire  sink_ACancel_earlyValid = idle ? _T_12 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [2:0] _GEN_21 = {{2'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [2:0] _beatsLeft_T_4 = beatsLeft - _GEN_21; // @[Arbiter.scala 113:52]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  out_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 123:31]
  wire [63:0] _T_29 = muxStateEarly_0 ? amo_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_30 = muxStateEarly_1 ? auto_in_a_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_32 = muxStateEarly_0 ? source_c_bits_a_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_33 = muxStateEarly_1 ? auto_in_a_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [30:0] _T_35 = muxStateEarly_0 ? cam_a_0_bits_address : 31'h0; // @[Mux.scala 27:73]
  wire [30:0] _T_36 = muxStateEarly_1 ? auto_in_a_bits_address : 31'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_38 = muxStateEarly_0 ? cam_a_0_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_39 = muxStateEarly_1 ? auto_in_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_41 = muxStateEarly_0 ? cam_a_0_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_42 = muxStateEarly_1 ? auto_in_a_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire  _T_50 = out_1_ready & source_i_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_39 = {{1'd0}, auto_in_a_bits_param[1:0]}; // @[Mux.scala 81:61]
  wire [3:0] _cam_a_0_lut_T_2 = 3'h1 == _GEN_39 ? 4'he : 4'h8; // @[Mux.scala 81:58]
  wire [1:0] _GEN_12 = cam_free_0 ? 2'h3 : cam_s_0_state; // @[AtomicAutomata.scala 187:23 188:23 76:28]
  wire [1:0] _GEN_23 = _T_50 & _T ? _GEN_12 : cam_s_0_state; // @[AtomicAutomata.scala 174:50 76:28]
  wire  _T_53 = out_ready & cam_amo_0; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_24 = cam_amo_0 ? 2'h1 : _GEN_23; // @[AtomicAutomata.scala 196:23 197:23]
  wire [1:0] _GEN_25 = _T_53 ? _GEN_24 : _GEN_23; // @[AtomicAutomata.scala 194:32]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25]
  wire  d_ackd = auto_out_d_bits_opcode == 3'h1; // @[AtomicAutomata.scala 213:40]
  wire  d_cam_sel_raw_0 = cam_a_0_bits_source == auto_out_d_bits_source; // @[AtomicAutomata.scala 204:53]
  wire  d_cam_sel_match_0 = d_cam_sel_raw_0 & cam_dmatch_0; // @[AtomicAutomata.scala 205:83]
  wire  d_drop = d_first & d_ackd & d_cam_sel_match_0; // @[AtomicAutomata.scala 232:40]
  wire  bundleOut_0_d_ready = auto_in_d_ready | d_drop; // @[AtomicAutomata.scala 236:35]
  wire  _d_first_T = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28]
  wire  d_ack = auto_out_d_bits_opcode == 3'h0; // @[AtomicAutomata.scala 214:40]
  wire  d_replace = d_first & d_ack & d_cam_sel_match_0; // @[AtomicAutomata.scala 233:42]
  reg [5:0] TLAtomicAutomata_covState; // @[Register tracking TLAtomicAutomata state]
  reg  TLAtomicAutomata_covMap [0:63]; // @[Coverage map for TLAtomicAutomata]
  wire  TLAtomicAutomata_covMap_read_en; // @[Coverage map for TLAtomicAutomata]
  wire [5:0] TLAtomicAutomata_covMap_read_addr; // @[Coverage map for TLAtomicAutomata]
  wire  TLAtomicAutomata_covMap_read_data; // @[Coverage map for TLAtomicAutomata]
  wire  TLAtomicAutomata_covMap_write_data; // @[Coverage map for TLAtomicAutomata]
  wire [5:0] TLAtomicAutomata_covMap_write_addr; // @[Coverage map for TLAtomicAutomata]
  wire  TLAtomicAutomata_covMap_write_mask; // @[Coverage map for TLAtomicAutomata]
  wire  TLAtomicAutomata_covMap_write_en; // @[Coverage map for TLAtomicAutomata]
  reg [29:0] TLAtomicAutomata_covSum; // @[Sum of coverage map]
  wire [1:0] cam_s_0_state_shl;
  wire [5:0] cam_s_0_state_pad;
  wire [4:0] d_first_counter_shl;
  wire [5:0] d_first_counter_pad;
  wire [5:0] state_0_shl;
  wire [5:0] state_0_pad;
  wire [5:0] state_1_shl;
  wire [5:0] state_1_pad;
  wire [5:0] TLAtomicAutomata_xor1;
  wire [5:0] TLAtomicAutomata_xor2;
  wire [5:0] TLAtomicAutomata_xor0;
  assign auto_in_a_ready = out_1_ready & a_allow; // @[AtomicAutomata.scala 150:38]
  assign auto_in_d_valid = auto_out_d_valid & ~d_drop; // @[AtomicAutomata.scala 235:35]
  assign auto_in_d_bits_opcode = d_replace ? 3'h1 : auto_out_d_bits_opcode; // @[AtomicAutomata.scala 238:19 239:26 240:28]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = d_replace ? cam_d_0_denied | auto_out_d_bits_denied : auto_out_d_bits_denied; // @[AtomicAutomata.scala 238:19 239:26 243:29]
  assign auto_in_d_bits_data = d_replace ? cam_d_0_data : auto_out_d_bits_data; // @[AtomicAutomata.scala 238:19 239:26 241:26]
  assign auto_in_d_bits_corrupt = d_replace ? cam_d_0_corrupt | auto_out_d_bits_denied : auto_out_d_bits_corrupt; // @[AtomicAutomata.scala 238:19 239:26 242:29]
  assign auto_out_a_valid = idle ? _T_12 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_out_a_bits_opcode = muxStateEarly_1 ? source_i_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  assign auto_out_a_bits_param = muxStateEarly_1 ? source_i_bits_param : 3'h0; // @[Mux.scala 27:73]
  assign auto_out_a_bits_size = _T_41 | _T_42; // @[Mux.scala 27:73]
  assign auto_out_a_bits_source = _T_38 | _T_39; // @[Mux.scala 27:73]
  assign auto_out_a_bits_address = _T_35 | _T_36; // @[Mux.scala 27:73]
  assign auto_out_a_bits_mask = _T_32 | _T_33; // @[Mux.scala 27:73]
  assign auto_out_a_bits_data = _T_29 | _T_30; // @[Mux.scala 27:73]
  assign auto_out_d_ready = auto_in_d_ready | d_drop; // @[AtomicAutomata.scala 236:35]
  assign TLAtomicAutomata_covMap_read_en = 1'h1;
  assign TLAtomicAutomata_covMap_read_addr = TLAtomicAutomata_covState;
  assign TLAtomicAutomata_covMap_read_data = TLAtomicAutomata_covMap[TLAtomicAutomata_covMap_read_addr]; // @[Coverage map for TLAtomicAutomata]
  assign TLAtomicAutomata_covMap_write_data = 1'h1;
  assign TLAtomicAutomata_covMap_write_addr = TLAtomicAutomata_covState;
  assign TLAtomicAutomata_covMap_write_mask = 1'h1;
  assign TLAtomicAutomata_covMap_write_en = ~metaReset;
  assign cam_s_0_state_shl = cam_s_0_state;
  assign cam_s_0_state_pad = {4'h0,cam_s_0_state_shl};
  assign d_first_counter_shl = {d_first_counter, 2'h0};
  assign d_first_counter_pad = {1'h0,d_first_counter_shl};
  assign state_0_shl = {state_0, 5'h0};
  assign state_0_pad = state_0_shl;
  assign state_1_shl = {state_1, 5'h0};
  assign state_1_pad = state_1_shl;
  assign TLAtomicAutomata_xor1 = cam_s_0_state_pad ^ d_first_counter_pad;
  assign TLAtomicAutomata_xor2 = state_0_pad ^ state_1_pad;
  assign TLAtomicAutomata_xor0 = TLAtomicAutomata_xor1 ^ TLAtomicAutomata_xor2;
  assign io_covSum = TLAtomicAutomata_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[AtomicAutomata.scala 76:28]
      cam_s_0_state <= 2'h0; // @[AtomicAutomata.scala 76:28]
    end else if (_d_first_T & d_first) begin
      if (d_cam_sel_match_0) begin
        if (d_ackd) begin
          cam_s_0_state <= 2'h2;
        end else begin
          cam_s_0_state <= 2'h0;
        end
      end else begin
        cam_s_0_state <= _GEN_25;
      end
    end else begin
      cam_s_0_state <= _GEN_25;
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_opcode <= auto_in_a_bits_opcode;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_param <= auto_in_a_bits_param;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_size <= auto_in_a_bits_size;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_source <= auto_in_a_bits_source;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_address <= auto_in_a_bits_address;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_mask <= auto_in_a_bits_mask;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_data <= auto_in_a_bits_data;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        if (3'h3 == _GEN_39) begin
          cam_a_0_lut <= 4'hc;
        end else if (3'h0 == _GEN_39) begin
          cam_a_0_lut <= 4'h6;
        end else begin
          cam_a_0_lut <= _cam_a_0_lut_T_2;
        end
      end
    end
    if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0 & d_ackd) begin
        cam_d_0_data <= auto_out_d_bits_data;
      end
    end
    if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0 & d_ackd) begin
        cam_d_0_denied <= auto_out_d_bits_denied;
      end
    end
    if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0 & d_ackd) begin
        cam_d_0_corrupt <= auto_out_d_bits_corrupt;
      end
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 3'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin
      if (earlyWinner_1) begin
        if (opdata) begin
          beatsLeft <= decode;
        end else begin
          beatsLeft <= 3'h0;
        end
      end else begin
        beatsLeft <= 3'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin
      if (d_first) begin
        if (d_first_beats1_opdata) begin
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1) & ~reset) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~earlyWinner_0 | ~earlyWinner_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(cam_amo_0 | source_i_valid) | (earlyWinner_0 | earlyWinner_1)) & _T_10) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(cam_amo_0 | source_i_valid) | (earlyWinner_0 | earlyWinner_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_13 | _T_12) & _T_10) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(_T_13 | _T_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    TLAtomicAutomata_covState <= TLAtomicAutomata_xor0;
    if (TLAtomicAutomata_covMap_write_en & TLAtomicAutomata_covMap_write_mask) begin
      TLAtomicAutomata_covMap[TLAtomicAutomata_covMap_write_addr] <= TLAtomicAutomata_covMap_write_data; // @[Coverage map for TLAtomicAutomata]
    end
    if (!(TLAtomicAutomata_covMap_read_data | metaReset)) begin
      TLAtomicAutomata_covSum <= TLAtomicAutomata_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    TLAtomicAutomata_covMap[initvar] = 0; //_17[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cam_s_0_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cam_a_0_bits_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  cam_a_0_bits_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  cam_a_0_bits_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  cam_a_0_bits_source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  cam_a_0_bits_address = _RAND_5[30:0];
  _RAND_6 = {1{`RANDOM}};
  cam_a_0_bits_mask = _RAND_6[7:0];
  _RAND_7 = {2{`RANDOM}};
  cam_a_0_bits_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  cam_a_0_lut = _RAND_8[3:0];
  _RAND_9 = {2{`RANDOM}};
  cam_d_0_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  cam_d_0_denied = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cam_d_0_corrupt = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  beatsLeft = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  state_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  d_first_counter = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  TLAtomicAutomata_covState = 0; //_16[5:0];
  _RAND_18 = {1{`RANDOM}};
  TLAtomicAutomata_covSum = 0; //_18[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [30:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [30:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [6:0] saved_source; // @[Repeater.scala 20:18]
  reg [30:0] saved_address; // @[Repeater.scala 20:18]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 19:21 28:{38,45}]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  reg  Repeater_covState; // @[Register tracking Repeater state]
  reg  Repeater_covMap [0:1]; // @[Coverage map for Repeater]
  wire  Repeater_covMap_read_en; // @[Coverage map for Repeater]
  wire  Repeater_covMap_read_addr; // @[Coverage map for Repeater]
  wire  Repeater_covMap_read_data; // @[Coverage map for Repeater]
  wire  Repeater_covMap_write_data; // @[Coverage map for Repeater]
  wire  Repeater_covMap_write_addr; // @[Coverage map for Repeater]
  wire  Repeater_covMap_write_mask; // @[Coverage map for Repeater]
  wire  Repeater_covMap_write_en; // @[Coverage map for Repeater]
  reg [29:0] Repeater_covSum; // @[Sum of coverage map]
  wire  full_shl;
  wire  full_pad;
  assign io_full = full; // @[Repeater.scala 26:11]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21]
  assign Repeater_covMap_read_en = 1'h1;
  assign Repeater_covMap_read_addr = Repeater_covState;
  assign Repeater_covMap_read_data = Repeater_covMap[Repeater_covMap_read_addr]; // @[Coverage map for Repeater]
  assign Repeater_covMap_write_data = 1'h1;
  assign Repeater_covMap_write_addr = Repeater_covState;
  assign Repeater_covMap_write_mask = 1'h1;
  assign Repeater_covMap_write_en = ~metaReset;
  assign full_shl = full;
  assign full_pad = full_shl;
  assign io_covSum = Repeater_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin
      full <= 1'h0;
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62]
    end
    Repeater_covState <= full_pad;
    if (Repeater_covMap_write_en & Repeater_covMap_write_mask) begin
      Repeater_covMap[Repeater_covMap_write_addr] <= Repeater_covMap_write_data; // @[Coverage map for Repeater]
    end
    if (!(Repeater_covMap_read_data | metaReset)) begin
      Repeater_covSum <= Repeater_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Repeater_covMap[initvar] = 0; //_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_source = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  saved_address = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  saved_mask = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  Repeater_covState = 0; //_6[0:0];
  _RAND_8 = {1{`RANDOM}};
  Repeater_covSum = 0; //_8[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [30:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [1:0]  auto_out_a_bits_size,
  output [10:0] auto_out_a_bits_source,
  output [30:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_size,
  input  [10:0] auto_out_d_bits_source,
  input  [63:0] auto_out_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  repeater_clock; // @[Fragmenter.scala 262:30]
  wire  repeater_reset; // @[Fragmenter.scala 262:30]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_opcode; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30]
  wire [30:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_opcode; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30]
  wire [30:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30]
  wire [29:0] repeater_io_covSum; // @[Fragmenter.scala 262:30]
  wire  repeater_metaReset; // @[Fragmenter.scala 262:30]
  reg [2:0] acknum; // @[Fragmenter.scala 189:29]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24]
  reg  dToggle; // @[Fragmenter.scala 191:30]
  wire [2:0] dFragnum = auto_out_d_bits_source[2:0]; // @[Fragmenter.scala 192:41]
  wire  dFirst = acknum == 3'h0; // @[Fragmenter.scala 193:29]
  wire  dLast = dFragnum == 3'h0; // @[Fragmenter.scala 194:30]
  wire [3:0] dsizeOH = 4'h1 << auto_out_d_bits_size; // @[OneHot.scala 64:12]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[package.scala 234:46]
  wire  dHasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  _T_5 = ~reset; // @[Fragmenter.scala 202:16]
  wire  ack_decrement = dHasData | dsizeOH[3]; // @[Fragmenter.scala 204:32]
  wire [5:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[Fragmenter.scala 206:47]
  wire [5:0] _GEN_7 = {{3'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69]
  wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69]
  wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0}; // @[package.scala 232:35]
  wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h1; // @[package.scala 232:40]
  wire [6:0] _dFirst_size_T_4 = {1'h0,_dFirst_size_T_1}; // @[Cat.scala 31:58]
  wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4; // @[package.scala 232:53]
  wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5; // @[package.scala 232:51]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4]; // @[OneHot.scala 30:18]
  wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_7 = |dFirst_size_hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28]
  wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo; // @[OneHot.scala 32:28]
  wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_9 = |dFirst_size_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] dFirst_size = {_dFirst_size_T_7,_dFirst_size_T_9,_dFirst_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  drop = ~dHasData & ~dLast; // @[Fragmenter.scala 222:30]
  wire  bundleOut_0_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35]
  wire  _T_7 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_9 = {{2'd0}, ack_decrement}; // @[Fragmenter.scala 209:55]
  wire [2:0] _acknum_T_1 = acknum - _GEN_9; // @[Fragmenter.scala 209:55]
  wire [2:0] aFrag = repeater_io_deq_bits_size > 3'h3 ? 3'h3 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[package.scala 234:77]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[package.scala 234:46]
  wire  aHasData = ~repeater_io_deq_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] gennum; // @[Fragmenter.scala 291:29]
  wire  aFirst = gennum == 3'h0; // @[Fragmenter.scala 292:29]
  wire [2:0] _old_gennum1_T_2 = gennum - 3'h1; // @[Fragmenter.scala 293:79]
  wire [2:0] old_gennum1 = aFirst ? aOrigOH1[5:3] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30]
  wire [2:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28]
  wire [2:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26]
  reg  aToggle_r; // @[Reg.scala 16:16]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  aToggle = ~_GEN_5; // @[Fragmenter.scala 297:23]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 50:35]
  wire  _repeater_io_repeat_T = ~aHasData; // @[Fragmenter.scala 302:31]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 3'h0}; // @[Fragmenter.scala 304:65]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88]
  wire [5:0] _GEN_10 = {{3'd0}, aFragOH1}; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h7; // @[Fragmenter.scala 304:111]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51]
  wire [30:0] _GEN_11 = {{25'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49]
  wire [7:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,aToggle}; // @[Cat.scala 31:58]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17]
  wire [29:0] TLFragmenter_covSum;
  wire [29:0] repeater_sum;
  Repeater repeater ( // @[Fragmenter.scala 262:30]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_opcode(repeater_io_enq_bits_opcode),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_opcode(repeater_io_deq_bits_opcode),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_covSum(repeater_io_covSum),
    .metaReset(repeater_metaReset)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 Fragmenter.scala 263:25]
  assign auto_in_d_valid = auto_out_d_valid & ~drop; // @[Fragmenter.scala 224:36]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32]
  assign auto_in_d_bits_source = auto_out_d_bits_source[10:4]; // @[Fragmenter.scala 226:47]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 Fragmenter.scala 306:25]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 31:58]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11; // @[Fragmenter.scala 304:49]
  assign auto_out_a_bits_mask = repeater_io_full ? 8'hff : auto_in_a_bits_mask; // @[Fragmenter.scala 313:31]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35]
  assign repeater_clock = clock;
  assign repeater_reset = reset;
  assign repeater_io_repeat = ~aHasData & new_gennum != 3'h0; // @[Fragmenter.scala 302:41]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign TLFragmenter_covSum = 30'h0;
  assign repeater_sum = TLFragmenter_covSum + repeater_io_covSum;
  assign io_covSum = repeater_sum;
  assign repeater_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29]
      acknum <= 3'h0; // @[Fragmenter.scala 189:29]
    end else if (_T_7) begin
      if (dFirst) begin
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29]
      if (dFirst) begin
        dOrig <= dFirst_size;
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30]
    end else if (_T_7) begin
      if (dFirst) begin
        dToggle <= auto_out_d_bits_source[3];
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29]
      gennum <= 3'h0; // @[Fragmenter.scala 291:29]
    end else if (_T_8) begin
      gennum <= new_gennum;
    end
    if (aFirst) begin // @[Reg.scala 17:18]
      aToggle_r <= dToggle; // @[Reg.scala 17:22]
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Fragmenter.scala 202:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~repeater_io_full | _repeater_io_repeat_T) & _T_5) begin
          $fatal; // @[Fragmenter.scala 309:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(~repeater_io_full | _repeater_io_repeat_T)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:309 assert (!repeater.io.full || !aHasData)\n"
            ); // @[Fragmenter.scala 309:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_9 | repeater_io_deq_bits_mask == 8'hff) & _T_5) begin
          $fatal; // @[Fragmenter.scala 312:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(_T_9 | repeater_io_deq_bits_mask == 8'hff)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLInterconnectCoupler_4(
  input         clock,
  input         reset,
  input         auto_control_xing_out_a_ready,
  output        auto_control_xing_out_a_valid,
  output [2:0]  auto_control_xing_out_a_bits_opcode,
  output [1:0]  auto_control_xing_out_a_bits_size,
  output [10:0] auto_control_xing_out_a_bits_source,
  output [30:0] auto_control_xing_out_a_bits_address,
  output [7:0]  auto_control_xing_out_a_bits_mask,
  output [63:0] auto_control_xing_out_a_bits_data,
  output        auto_control_xing_out_d_ready,
  input         auto_control_xing_out_d_valid,
  input  [2:0]  auto_control_xing_out_d_bits_opcode,
  input  [1:0]  auto_control_xing_out_d_bits_size,
  input  [10:0] auto_control_xing_out_d_bits_source,
  input  [63:0] auto_control_xing_out_d_bits_data,
  output        auto_tl_in_a_ready,
  input         auto_tl_in_a_valid,
  input  [2:0]  auto_tl_in_a_bits_opcode,
  input  [2:0]  auto_tl_in_a_bits_size,
  input  [6:0]  auto_tl_in_a_bits_source,
  input  [30:0] auto_tl_in_a_bits_address,
  input  [7:0]  auto_tl_in_a_bits_mask,
  input  [63:0] auto_tl_in_a_bits_data,
  input         auto_tl_in_d_ready,
  output        auto_tl_in_d_valid,
  output [2:0]  auto_tl_in_d_bits_opcode,
  output [2:0]  auto_tl_in_d_bits_size,
  output [6:0]  auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [30:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_in_a_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_out_a_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [30:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [7:0] fragmenter_auto_out_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_out_a_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_out_d_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34]
  wire [29:0] fragmenter_io_covSum; // @[Fragmenter.scala 333:34]
  wire  fragmenter_metaReset; // @[Fragmenter.scala 333:34]
  wire [29:0] TLInterconnectCoupler_4_covSum;
  wire [29:0] fragmenter_sum;
  TLFragmenter fragmenter ( // @[Fragmenter.scala 333:34]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .io_covSum(fragmenter_io_covSum),
    .metaReset(fragmenter_metaReset)
  );
  assign auto_control_xing_out_a_valid = fragmenter_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_control_xing_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_control_xing_out_a_bits_size = fragmenter_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_control_xing_out_a_bits_source = fragmenter_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_control_xing_out_a_bits_address = fragmenter_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_control_xing_out_a_bits_mask = fragmenter_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_control_xing_out_a_bits_data = fragmenter_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_control_xing_out_d_ready = fragmenter_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_opcode = fragmenter_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign fragmenter_clock = clock;
  assign fragmenter_reset = reset;
  assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_data = auto_tl_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_out_a_ready = auto_control_xing_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_valid = auto_control_xing_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_opcode = auto_control_xing_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_size = auto_control_xing_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_source = auto_control_xing_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_data = auto_control_xing_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign TLInterconnectCoupler_4_covSum = 30'h0;
  assign fragmenter_sum = TLInterconnectCoupler_4_covSum + fragmenter_io_covSum;
  assign io_covSum = fragmenter_sum;
  assign fragmenter_metaReset = metaReset;
endmodule
module PeripheryBus(
  input         auto_coupler_to_device_named_uart_0_control_xing_out_a_ready,
  output        auto_coupler_to_device_named_uart_0_control_xing_out_a_valid,
  output [2:0]  auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode,
  output [1:0]  auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size,
  output [10:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source,
  output [30:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address,
  output [7:0]  auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask,
  output [63:0] auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data,
  output        auto_coupler_to_device_named_uart_0_control_xing_out_d_ready,
  input         auto_coupler_to_device_named_uart_0_control_xing_out_d_valid,
  input  [2:0]  auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode,
  input  [1:0]  auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size,
  input  [10:0] auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source,
  input  [63:0] auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data,
  output        auto_fixedClockNode_out_clock,
  output        auto_fixedClockNode_out_reset,
  input         auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock,
  input         auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset,
  output        auto_bus_xing_in_a_ready,
  input         auto_bus_xing_in_a_valid,
  input  [2:0]  auto_bus_xing_in_a_bits_opcode,
  input  [2:0]  auto_bus_xing_in_a_bits_param,
  input  [2:0]  auto_bus_xing_in_a_bits_size,
  input  [6:0]  auto_bus_xing_in_a_bits_source,
  input  [30:0] auto_bus_xing_in_a_bits_address,
  input  [7:0]  auto_bus_xing_in_a_bits_mask,
  input  [63:0] auto_bus_xing_in_a_bits_data,
  input         auto_bus_xing_in_d_ready,
  output        auto_bus_xing_in_d_valid,
  output [2:0]  auto_bus_xing_in_d_bits_opcode,
  output [2:0]  auto_bus_xing_in_d_bits_size,
  output [6:0]  auto_bus_xing_in_d_bits_source,
  output        auto_bus_xing_in_d_bits_denied,
  output [63:0] auto_bus_xing_in_d_bits_data,
  output        auto_bus_xing_in_d_bits_corrupt,
  output        clock,
  output        reset,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_clock;
  wire  subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_reset;
  wire  subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_clock;
  wire  subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_reset;
  wire  clockGroup_auto_in_member_subsystem_pbus_0_clock;
  wire  clockGroup_auto_in_member_subsystem_pbus_0_reset;
  wire  clockGroup_auto_out_clock;
  wire  clockGroup_auto_out_reset;
  wire  fixedClockNode_auto_in_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_in_reset; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_1_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_1_reset; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_0_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_0_reset; // @[ClockGroup.scala 106:107]
  wire [29:0] fixedClockNode_io_covSum; // @[ClockGroup.scala 106:107]
  wire  fixer_auto_in_a_ready; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_in_a_valid; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_in_a_bits_opcode; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_in_a_bits_size; // @[PeripheryBus.scala 47:33]
  wire [6:0] fixer_auto_in_a_bits_source; // @[PeripheryBus.scala 47:33]
  wire [30:0] fixer_auto_in_a_bits_address; // @[PeripheryBus.scala 47:33]
  wire [7:0] fixer_auto_in_a_bits_mask; // @[PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_in_a_bits_data; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_in_d_ready; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_in_d_valid; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_in_d_bits_opcode; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_in_d_bits_size; // @[PeripheryBus.scala 47:33]
  wire [6:0] fixer_auto_in_d_bits_source; // @[PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_in_d_bits_data; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_a_ready; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_a_valid; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_out_a_bits_opcode; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_out_a_bits_size; // @[PeripheryBus.scala 47:33]
  wire [6:0] fixer_auto_out_a_bits_source; // @[PeripheryBus.scala 47:33]
  wire [30:0] fixer_auto_out_a_bits_address; // @[PeripheryBus.scala 47:33]
  wire [7:0] fixer_auto_out_a_bits_mask; // @[PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_out_a_bits_data; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_d_ready; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_d_valid; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_out_d_bits_opcode; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_out_d_bits_size; // @[PeripheryBus.scala 47:33]
  wire [6:0] fixer_auto_out_d_bits_source; // @[PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_out_d_bits_data; // @[PeripheryBus.scala 47:33]
  wire [29:0] fixer_io_covSum; // @[PeripheryBus.scala 47:33]
  wire  in_xbar_auto_in_a_ready;
  wire  in_xbar_auto_in_a_valid;
  wire [2:0] in_xbar_auto_in_a_bits_opcode;
  wire [2:0] in_xbar_auto_in_a_bits_param;
  wire [2:0] in_xbar_auto_in_a_bits_size;
  wire [6:0] in_xbar_auto_in_a_bits_source;
  wire [30:0] in_xbar_auto_in_a_bits_address;
  wire [7:0] in_xbar_auto_in_a_bits_mask;
  wire [63:0] in_xbar_auto_in_a_bits_data;
  wire  in_xbar_auto_in_d_ready;
  wire  in_xbar_auto_in_d_valid;
  wire [2:0] in_xbar_auto_in_d_bits_opcode;
  wire [2:0] in_xbar_auto_in_d_bits_size;
  wire [6:0] in_xbar_auto_in_d_bits_source;
  wire  in_xbar_auto_in_d_bits_denied;
  wire [63:0] in_xbar_auto_in_d_bits_data;
  wire  in_xbar_auto_in_d_bits_corrupt;
  wire  in_xbar_auto_out_a_ready;
  wire  in_xbar_auto_out_a_valid;
  wire [2:0] in_xbar_auto_out_a_bits_opcode;
  wire [2:0] in_xbar_auto_out_a_bits_param;
  wire [2:0] in_xbar_auto_out_a_bits_size;
  wire [6:0] in_xbar_auto_out_a_bits_source;
  wire [30:0] in_xbar_auto_out_a_bits_address;
  wire [7:0] in_xbar_auto_out_a_bits_mask;
  wire [63:0] in_xbar_auto_out_a_bits_data;
  wire  in_xbar_auto_out_d_ready;
  wire  in_xbar_auto_out_d_valid;
  wire [2:0] in_xbar_auto_out_d_bits_opcode;
  wire [2:0] in_xbar_auto_out_d_bits_size;
  wire [6:0] in_xbar_auto_out_d_bits_source;
  wire  in_xbar_auto_out_d_bits_denied;
  wire [63:0] in_xbar_auto_out_d_bits_data;
  wire  in_xbar_auto_out_d_bits_corrupt;
  wire  out_xbar_auto_in_a_ready;
  wire  out_xbar_auto_in_a_valid;
  wire [2:0] out_xbar_auto_in_a_bits_opcode;
  wire [2:0] out_xbar_auto_in_a_bits_size;
  wire [6:0] out_xbar_auto_in_a_bits_source;
  wire [30:0] out_xbar_auto_in_a_bits_address;
  wire [7:0] out_xbar_auto_in_a_bits_mask;
  wire [63:0] out_xbar_auto_in_a_bits_data;
  wire  out_xbar_auto_in_d_ready;
  wire  out_xbar_auto_in_d_valid;
  wire [2:0] out_xbar_auto_in_d_bits_opcode;
  wire [2:0] out_xbar_auto_in_d_bits_size;
  wire [6:0] out_xbar_auto_in_d_bits_source;
  wire [63:0] out_xbar_auto_in_d_bits_data;
  wire  out_xbar_auto_out_a_ready;
  wire  out_xbar_auto_out_a_valid;
  wire [2:0] out_xbar_auto_out_a_bits_opcode;
  wire [2:0] out_xbar_auto_out_a_bits_size;
  wire [6:0] out_xbar_auto_out_a_bits_source;
  wire [30:0] out_xbar_auto_out_a_bits_address;
  wire [7:0] out_xbar_auto_out_a_bits_mask;
  wire [63:0] out_xbar_auto_out_a_bits_data;
  wire  out_xbar_auto_out_d_ready;
  wire  out_xbar_auto_out_d_valid;
  wire [2:0] out_xbar_auto_out_d_bits_opcode;
  wire [2:0] out_xbar_auto_out_d_bits_size;
  wire [6:0] out_xbar_auto_out_d_bits_source;
  wire [63:0] out_xbar_auto_out_d_bits_data;
  wire  buffer_clock; // @[Buffer.scala 68:28]
  wire  buffer_reset; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28]
  wire [30:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28]
  wire [30:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire [29:0] buffer_io_covSum; // @[Buffer.scala 68:28]
  wire  atomics_clock; // @[AtomicAutomata.scala 283:29]
  wire  atomics_reset; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_a_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_a_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_a_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_a_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_a_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_in_a_bits_source; // @[AtomicAutomata.scala 283:29]
  wire [30:0] atomics_auto_in_a_bits_address; // @[AtomicAutomata.scala 283:29]
  wire [7:0] atomics_auto_in_a_bits_mask; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_in_a_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_d_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_d_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_in_d_bits_source; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_bits_denied; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_in_d_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_bits_corrupt; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_a_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_a_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_a_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_a_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_a_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_out_a_bits_source; // @[AtomicAutomata.scala 283:29]
  wire [30:0] atomics_auto_out_a_bits_address; // @[AtomicAutomata.scala 283:29]
  wire [7:0] atomics_auto_out_a_bits_mask; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_out_a_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_d_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_d_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_out_d_bits_source; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_bits_denied; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_out_d_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_bits_corrupt; // @[AtomicAutomata.scala 283:29]
  wire [29:0] atomics_io_covSum; // @[AtomicAutomata.scala 283:29]
  wire  atomics_metaReset; // @[AtomicAutomata.scala 283:29]
  wire  buffer_1_clock; // @[Buffer.scala 68:28]
  wire  buffer_1_reset; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_in_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_in_a_bits_param; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_in_a_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_1_auto_in_a_bits_source; // @[Buffer.scala 68:28]
  wire [30:0] buffer_1_auto_in_a_bits_address; // @[Buffer.scala 68:28]
  wire [7:0] buffer_1_auto_in_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_1_auto_in_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_in_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_in_d_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_1_auto_in_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_1_auto_in_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_out_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_out_a_bits_param; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_out_a_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_1_auto_out_a_bits_source; // @[Buffer.scala 68:28]
  wire [30:0] buffer_1_auto_out_a_bits_address; // @[Buffer.scala 68:28]
  wire [7:0] buffer_1_auto_out_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_1_auto_out_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_out_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_out_d_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_1_auto_out_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_1_auto_out_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire [29:0] buffer_1_io_covSum; // @[Buffer.scala 68:28]
  wire  coupler_to_device_named_uart_0_clock; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_reset; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_auto_control_xing_out_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_auto_control_xing_out_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_source; // @[LazyModule.scala 432:27]
  wire [30:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_mask; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_auto_control_xing_out_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_auto_control_xing_out_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_auto_tl_in_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_auto_tl_in_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_source; // @[LazyModule.scala 432:27]
  wire [30:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_mask; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_device_named_uart_0_auto_tl_in_a_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_auto_tl_in_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_auto_tl_in_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_device_named_uart_0_auto_tl_in_d_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_device_named_uart_0_auto_tl_in_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_device_named_uart_0_auto_tl_in_d_bits_data; // @[LazyModule.scala 432:27]
  wire [29:0] coupler_to_device_named_uart_0_io_covSum; // @[LazyModule.scala 432:27]
  wire  coupler_to_device_named_uart_0_metaReset; // @[LazyModule.scala 432:27]
  wire [29:0] PeripheryBus_covSum;
  wire [29:0] buffer_sum;
  wire [29:0] fixedClockNode_sum;
  wire [29:0] fixer_sum;
  wire [29:0] buffer_1_sum;
  wire [29:0] coupler_to_device_named_uart_0_sum;
  wire [29:0] atomics_sum;
  FixedClockBroadcast_1 fixedClockNode ( // @[ClockGroup.scala 106:107]
    .auto_in_clock(fixedClockNode_auto_in_clock),
    .auto_in_reset(fixedClockNode_auto_in_reset),
    .auto_out_1_clock(fixedClockNode_auto_out_1_clock),
    .auto_out_1_reset(fixedClockNode_auto_out_1_reset),
    .auto_out_0_clock(fixedClockNode_auto_out_0_clock),
    .auto_out_0_reset(fixedClockNode_auto_out_0_reset),
    .io_covSum(fixedClockNode_io_covSum)
  );
  TLFIFOFixer_1 fixer ( // @[PeripheryBus.scala 47:33]
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_auto_in_a_bits_data),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_auto_out_a_bits_data),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data),
    .io_covSum(fixer_io_covSum)
  );
  TLBuffer buffer ( // @[Buffer.scala 68:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt),
    .io_covSum(buffer_io_covSum)
  );
  TLAtomicAutomata atomics ( // @[AtomicAutomata.scala 283:29]
    .clock(atomics_clock),
    .reset(atomics_reset),
    .auto_in_a_ready(atomics_auto_in_a_ready),
    .auto_in_a_valid(atomics_auto_in_a_valid),
    .auto_in_a_bits_opcode(atomics_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(atomics_auto_in_a_bits_param),
    .auto_in_a_bits_size(atomics_auto_in_a_bits_size),
    .auto_in_a_bits_source(atomics_auto_in_a_bits_source),
    .auto_in_a_bits_address(atomics_auto_in_a_bits_address),
    .auto_in_a_bits_mask(atomics_auto_in_a_bits_mask),
    .auto_in_a_bits_data(atomics_auto_in_a_bits_data),
    .auto_in_d_ready(atomics_auto_in_d_ready),
    .auto_in_d_valid(atomics_auto_in_d_valid),
    .auto_in_d_bits_opcode(atomics_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(atomics_auto_in_d_bits_size),
    .auto_in_d_bits_source(atomics_auto_in_d_bits_source),
    .auto_in_d_bits_denied(atomics_auto_in_d_bits_denied),
    .auto_in_d_bits_data(atomics_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(atomics_auto_in_d_bits_corrupt),
    .auto_out_a_ready(atomics_auto_out_a_ready),
    .auto_out_a_valid(atomics_auto_out_a_valid),
    .auto_out_a_bits_opcode(atomics_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(atomics_auto_out_a_bits_param),
    .auto_out_a_bits_size(atomics_auto_out_a_bits_size),
    .auto_out_a_bits_source(atomics_auto_out_a_bits_source),
    .auto_out_a_bits_address(atomics_auto_out_a_bits_address),
    .auto_out_a_bits_mask(atomics_auto_out_a_bits_mask),
    .auto_out_a_bits_data(atomics_auto_out_a_bits_data),
    .auto_out_d_ready(atomics_auto_out_d_ready),
    .auto_out_d_valid(atomics_auto_out_d_valid),
    .auto_out_d_bits_opcode(atomics_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(atomics_auto_out_d_bits_size),
    .auto_out_d_bits_source(atomics_auto_out_d_bits_source),
    .auto_out_d_bits_denied(atomics_auto_out_d_bits_denied),
    .auto_out_d_bits_data(atomics_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(atomics_auto_out_d_bits_corrupt),
    .io_covSum(atomics_io_covSum),
    .metaReset(atomics_metaReset)
  );
  TLBuffer buffer_1 ( // @[Buffer.scala 68:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_a_ready(buffer_1_auto_in_a_ready),
    .auto_in_a_valid(buffer_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_1_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_1_auto_in_d_ready),
    .auto_in_d_valid(buffer_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(buffer_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_1_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_1_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_1_auto_out_a_ready),
    .auto_out_a_valid(buffer_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
    .auto_out_d_ready(buffer_1_auto_out_d_ready),
    .auto_out_d_valid(buffer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
    .auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt),
    .io_covSum(buffer_1_io_covSum)
  );
  TLInterconnectCoupler_4 coupler_to_device_named_uart_0 ( // @[LazyModule.scala 432:27]
    .clock(coupler_to_device_named_uart_0_clock),
    .reset(coupler_to_device_named_uart_0_reset),
    .auto_control_xing_out_a_ready(coupler_to_device_named_uart_0_auto_control_xing_out_a_ready),
    .auto_control_xing_out_a_valid(coupler_to_device_named_uart_0_auto_control_xing_out_a_valid),
    .auto_control_xing_out_a_bits_opcode(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_opcode),
    .auto_control_xing_out_a_bits_size(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_size),
    .auto_control_xing_out_a_bits_source(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_source),
    .auto_control_xing_out_a_bits_address(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_address),
    .auto_control_xing_out_a_bits_mask(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_mask),
    .auto_control_xing_out_a_bits_data(coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_data),
    .auto_control_xing_out_d_ready(coupler_to_device_named_uart_0_auto_control_xing_out_d_ready),
    .auto_control_xing_out_d_valid(coupler_to_device_named_uart_0_auto_control_xing_out_d_valid),
    .auto_control_xing_out_d_bits_opcode(coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_opcode),
    .auto_control_xing_out_d_bits_size(coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_size),
    .auto_control_xing_out_d_bits_source(coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_source),
    .auto_control_xing_out_d_bits_data(coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_data),
    .auto_tl_in_a_ready(coupler_to_device_named_uart_0_auto_tl_in_a_ready),
    .auto_tl_in_a_valid(coupler_to_device_named_uart_0_auto_tl_in_a_valid),
    .auto_tl_in_a_bits_opcode(coupler_to_device_named_uart_0_auto_tl_in_a_bits_opcode),
    .auto_tl_in_a_bits_size(coupler_to_device_named_uart_0_auto_tl_in_a_bits_size),
    .auto_tl_in_a_bits_source(coupler_to_device_named_uart_0_auto_tl_in_a_bits_source),
    .auto_tl_in_a_bits_address(coupler_to_device_named_uart_0_auto_tl_in_a_bits_address),
    .auto_tl_in_a_bits_mask(coupler_to_device_named_uart_0_auto_tl_in_a_bits_mask),
    .auto_tl_in_a_bits_data(coupler_to_device_named_uart_0_auto_tl_in_a_bits_data),
    .auto_tl_in_d_ready(coupler_to_device_named_uart_0_auto_tl_in_d_ready),
    .auto_tl_in_d_valid(coupler_to_device_named_uart_0_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_opcode(coupler_to_device_named_uart_0_auto_tl_in_d_bits_opcode),
    .auto_tl_in_d_bits_size(coupler_to_device_named_uart_0_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source(coupler_to_device_named_uart_0_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_data(coupler_to_device_named_uart_0_auto_tl_in_d_bits_data),
    .io_covSum(coupler_to_device_named_uart_0_io_covSum),
    .metaReset(coupler_to_device_named_uart_0_metaReset)
  );
  assign subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_clock =
    subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_reset =
    subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_clock = clockGroup_auto_in_member_subsystem_pbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_reset = clockGroup_auto_in_member_subsystem_pbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_in_a_ready = in_xbar_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_valid = in_xbar_auto_out_d_valid; // @[ReadyValidCancel.scala 21:38]
  assign in_xbar_auto_in_d_bits_opcode = in_xbar_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_bits_size = in_xbar_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_bits_source = in_xbar_auto_out_d_bits_source; // @[Xbar.scala 228:69]
  assign in_xbar_auto_in_d_bits_denied = in_xbar_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_bits_data = in_xbar_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_bits_corrupt = in_xbar_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_out_a_valid = in_xbar_auto_in_a_valid; // @[ReadyValidCancel.scala 21:38]
  assign in_xbar_auto_out_a_bits_opcode = in_xbar_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_param = in_xbar_auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_size = in_xbar_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_source = in_xbar_auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign in_xbar_auto_out_a_bits_address = in_xbar_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_mask = in_xbar_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_data = in_xbar_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_d_ready = in_xbar_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_xbar_auto_in_a_ready = out_xbar_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign out_xbar_auto_in_d_valid = out_xbar_auto_out_d_valid; // @[ReadyValidCancel.scala 21:38]
  assign out_xbar_auto_in_d_bits_opcode = out_xbar_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign out_xbar_auto_in_d_bits_size = out_xbar_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign out_xbar_auto_in_d_bits_source = out_xbar_auto_out_d_bits_source; // @[Xbar.scala 228:69]
  assign out_xbar_auto_in_d_bits_data = out_xbar_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign out_xbar_auto_out_a_valid = out_xbar_auto_in_a_valid; // @[ReadyValidCancel.scala 21:38]
  assign out_xbar_auto_out_a_bits_opcode = out_xbar_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_xbar_auto_out_a_bits_size = out_xbar_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_xbar_auto_out_a_bits_source = out_xbar_auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign out_xbar_auto_out_a_bits_address = out_xbar_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_xbar_auto_out_a_bits_mask = out_xbar_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_xbar_auto_out_a_bits_data = out_xbar_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_xbar_auto_out_d_ready = out_xbar_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_coupler_to_device_named_uart_0_control_xing_out_a_valid =
    coupler_to_device_named_uart_0_auto_control_xing_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode =
    coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size =
    coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source =
    coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address =
    coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask =
    coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data =
    coupler_to_device_named_uart_0_auto_control_xing_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_device_named_uart_0_control_xing_out_d_ready =
    coupler_to_device_named_uart_0_auto_control_xing_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_fixedClockNode_out_clock = fixedClockNode_auto_out_1_clock; // @[LazyModule.scala 311:12]
  assign auto_fixedClockNode_out_reset = fixedClockNode_auto_out_1_reset; // @[LazyModule.scala 311:12]
  assign auto_bus_xing_in_a_ready = buffer_1_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_valid = buffer_1_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_opcode = buffer_1_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_size = buffer_1_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_source = buffer_1_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_denied = buffer_1_auto_in_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_data = buffer_1_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_corrupt = buffer_1_auto_in_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_clock =
    auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock; // @[LazyModule.scala 309:16]
  assign subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_reset =
    auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset; // @[LazyModule.scala 309:16]
  assign clockGroup_auto_in_member_subsystem_pbus_0_clock =
    subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_clock; // @[LazyModule.scala 298:16]
  assign clockGroup_auto_in_member_subsystem_pbus_0_reset =
    subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_reset; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[LazyModule.scala 298:16]
  assign fixer_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_a_ready = out_xbar_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_valid = out_xbar_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_opcode = out_xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_size = out_xbar_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_source = out_xbar_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_data = out_xbar_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_in_a_valid = buffer_1_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_param = buffer_1_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_size = buffer_1_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_source = buffer_1_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_address = buffer_1_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_mask = buffer_1_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_data = buffer_1_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_d_ready = buffer_1_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_out_a_ready = atomics_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_valid = atomics_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_opcode = atomics_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_size = atomics_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_source = atomics_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_denied = atomics_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_data = atomics_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_corrupt = atomics_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_valid = fixer_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_size = fixer_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_source = fixer_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_address = fixer_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_data = fixer_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_d_ready = fixer_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_a_ready = coupler_to_device_named_uart_0_auto_tl_in_a_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_d_valid = coupler_to_device_named_uart_0_auto_tl_in_d_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_d_bits_opcode = coupler_to_device_named_uart_0_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_d_bits_size = coupler_to_device_named_uart_0_auto_tl_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_d_bits_source = coupler_to_device_named_uart_0_auto_tl_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_d_bits_data = coupler_to_device_named_uart_0_auto_tl_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign buffer_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign buffer_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign buffer_auto_in_a_valid = atomics_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_opcode = atomics_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_param = atomics_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_size = atomics_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_source = atomics_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_address = atomics_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_mask = atomics_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_data = atomics_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_d_ready = atomics_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_a_ready = fixer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_valid = fixer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_size = fixer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_source = fixer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_denied = 1'h0; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_data = fixer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_corrupt = 1'h0; // @[LazyModule.scala 296:16]
  assign atomics_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign atomics_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign atomics_auto_in_a_valid = in_xbar_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_opcode = in_xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_param = in_xbar_auto_out_a_bits_param; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_size = in_xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_source = in_xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_address = in_xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_mask = in_xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_data = in_xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_d_ready = in_xbar_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign atomics_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign buffer_1_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign buffer_1_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign buffer_1_auto_in_a_valid = auto_bus_xing_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_opcode = auto_bus_xing_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_param = auto_bus_xing_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_size = auto_bus_xing_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_source = auto_bus_xing_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_address = auto_bus_xing_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_mask = auto_bus_xing_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_data = auto_bus_xing_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_d_ready = auto_bus_xing_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_a_ready = in_xbar_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_valid = in_xbar_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_opcode = in_xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_size = in_xbar_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_source = in_xbar_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_denied = in_xbar_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_data = in_xbar_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_corrupt = in_xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign coupler_to_device_named_uart_0_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_device_named_uart_0_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_device_named_uart_0_auto_control_xing_out_a_ready =
    auto_coupler_to_device_named_uart_0_control_xing_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_device_named_uart_0_auto_control_xing_out_d_valid =
    auto_coupler_to_device_named_uart_0_control_xing_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_opcode =
    auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_size =
    auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_source =
    auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_device_named_uart_0_auto_control_xing_out_d_bits_data =
    auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_device_named_uart_0_auto_tl_in_a_valid = out_xbar_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_opcode = out_xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_size = out_xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_source = out_xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_address = out_xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_mask = out_xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_device_named_uart_0_auto_tl_in_a_bits_data = out_xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign coupler_to_device_named_uart_0_auto_tl_in_d_ready = out_xbar_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign PeripheryBus_covSum = 30'h0;
  assign buffer_sum = PeripheryBus_covSum + buffer_io_covSum;
  assign fixedClockNode_sum = buffer_sum + fixedClockNode_io_covSum;
  assign fixer_sum = fixedClockNode_sum + fixer_io_covSum;
  assign buffer_1_sum = fixer_sum + buffer_1_io_covSum;
  assign coupler_to_device_named_uart_0_sum = buffer_1_sum + coupler_to_device_named_uart_0_io_covSum;
  assign atomics_sum = coupler_to_device_named_uart_0_sum + atomics_io_covSum;
  assign io_covSum = atomics_sum;
  assign coupler_to_device_named_uart_0_metaReset = metaReset;
  assign atomics_metaReset = metaReset;
endmodule
module Queue_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input         io_enq_bits_user_amba_prot_bufferable,
  input         io_enq_bits_user_amba_prot_modifiable,
  input         io_enq_bits_user_amba_prot_readalloc,
  input         io_enq_bits_user_amba_prot_writealloc,
  input         io_enq_bits_user_amba_prot_privileged,
  input         io_enq_bits_user_amba_prot_secure,
  input         io_enq_bits_user_amba_prot_fetch,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output        io_deq_bits_user_amba_prot_bufferable,
  output        io_deq_bits_user_amba_prot_modifiable,
  output        io_deq_bits_user_amba_prot_readalloc,
  output        io_deq_bits_user_amba_prot_writealloc,
  output        io_deq_bits_user_amba_prot_privileged,
  output        io_deq_bits_user_amba_prot_secure,
  output        io_deq_bits_user_amba_prot_fetch,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_param_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_bufferable [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_modifiable [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_readalloc [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_writealloc [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_privileged [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_secure [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_fetch [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_4_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_en = 1'h1;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_bufferable_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_bufferable_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_bufferable_io_deq_bits_MPORT_data =
    ram_user_amba_prot_bufferable[ram_user_amba_prot_bufferable_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_bufferable_MPORT_data = io_enq_bits_user_amba_prot_bufferable;
  assign ram_user_amba_prot_bufferable_MPORT_addr = value;
  assign ram_user_amba_prot_bufferable_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_bufferable_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_modifiable_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_modifiable_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_modifiable_io_deq_bits_MPORT_data =
    ram_user_amba_prot_modifiable[ram_user_amba_prot_modifiable_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_modifiable_MPORT_data = io_enq_bits_user_amba_prot_modifiable;
  assign ram_user_amba_prot_modifiable_MPORT_addr = value;
  assign ram_user_amba_prot_modifiable_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_modifiable_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_readalloc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_readalloc_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_readalloc_io_deq_bits_MPORT_data =
    ram_user_amba_prot_readalloc[ram_user_amba_prot_readalloc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_readalloc_MPORT_data = io_enq_bits_user_amba_prot_readalloc;
  assign ram_user_amba_prot_readalloc_MPORT_addr = value;
  assign ram_user_amba_prot_readalloc_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_readalloc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_writealloc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_writealloc_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_writealloc_io_deq_bits_MPORT_data =
    ram_user_amba_prot_writealloc[ram_user_amba_prot_writealloc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_writealloc_MPORT_data = io_enq_bits_user_amba_prot_writealloc;
  assign ram_user_amba_prot_writealloc_MPORT_addr = value;
  assign ram_user_amba_prot_writealloc_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_writealloc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_privileged_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_privileged_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_privileged_io_deq_bits_MPORT_data =
    ram_user_amba_prot_privileged[ram_user_amba_prot_privileged_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_privileged_MPORT_data = io_enq_bits_user_amba_prot_privileged;
  assign ram_user_amba_prot_privileged_MPORT_addr = value;
  assign ram_user_amba_prot_privileged_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_privileged_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_secure_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_secure_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_secure_io_deq_bits_MPORT_data =
    ram_user_amba_prot_secure[ram_user_amba_prot_secure_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_secure_MPORT_data = io_enq_bits_user_amba_prot_secure;
  assign ram_user_amba_prot_secure_MPORT_addr = value;
  assign ram_user_amba_prot_secure_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_secure_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_fetch_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_fetch_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_fetch_io_deq_bits_MPORT_data =
    ram_user_amba_prot_fetch[ram_user_amba_prot_fetch_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_fetch_MPORT_data = io_enq_bits_user_amba_prot_fetch;
  assign ram_user_amba_prot_fetch_MPORT_addr = value;
  assign ram_user_amba_prot_fetch_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_fetch_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_bufferable = ram_user_amba_prot_bufferable_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_modifiable = ram_user_amba_prot_modifiable_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_readalloc = ram_user_amba_prot_readalloc_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_writealloc = ram_user_amba_prot_writealloc_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_privileged = ram_user_amba_prot_privileged_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_secure = ram_user_amba_prot_secure_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_fetch = ram_user_amba_prot_fetch_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_4_covSum = 30'h0;
  assign io_covSum = Queue_4_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_bufferable_MPORT_en & ram_user_amba_prot_bufferable_MPORT_mask) begin
      ram_user_amba_prot_bufferable[ram_user_amba_prot_bufferable_MPORT_addr] <=
        ram_user_amba_prot_bufferable_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_modifiable_MPORT_en & ram_user_amba_prot_modifiable_MPORT_mask) begin
      ram_user_amba_prot_modifiable[ram_user_amba_prot_modifiable_MPORT_addr] <=
        ram_user_amba_prot_modifiable_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_readalloc_MPORT_en & ram_user_amba_prot_readalloc_MPORT_mask) begin
      ram_user_amba_prot_readalloc[ram_user_amba_prot_readalloc_MPORT_addr] <= ram_user_amba_prot_readalloc_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_writealloc_MPORT_en & ram_user_amba_prot_writealloc_MPORT_mask) begin
      ram_user_amba_prot_writealloc[ram_user_amba_prot_writealloc_MPORT_addr] <=
        ram_user_amba_prot_writealloc_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_privileged_MPORT_en & ram_user_amba_prot_privileged_MPORT_mask) begin
      ram_user_amba_prot_privileged[ram_user_amba_prot_privileged_MPORT_addr] <=
        ram_user_amba_prot_privileged_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_secure_MPORT_en & ram_user_amba_prot_secure_MPORT_mask) begin
      ram_user_amba_prot_secure[ram_user_amba_prot_secure_MPORT_addr] <= ram_user_amba_prot_secure_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_fetch_MPORT_en & ram_user_amba_prot_fetch_MPORT_mask) begin
      ram_user_amba_prot_fetch[ram_user_amba_prot_fetch_MPORT_addr] <= ram_user_amba_prot_fetch_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= value_1 + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_bufferable[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_modifiable[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_readalloc[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_writealloc[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_privileged[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_secure[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_fetch[initvar] = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_12[7:0];
  _RAND_13 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_13[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  value = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  value_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  maybe_full = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_5(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [3:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input         io_enq_bits_denied,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [3:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output        io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_denied [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_5_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_5_covSum = 30'h0;
  assign io_covSum = Queue_5_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= value_1 + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_5[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  value_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_2(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [3:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input         auto_in_a_bits_user_amba_prot_bufferable,
  input         auto_in_a_bits_user_amba_prot_modifiable,
  input         auto_in_a_bits_user_amba_prot_readalloc,
  input         auto_in_a_bits_user_amba_prot_writealloc,
  input         auto_in_a_bits_user_amba_prot_privileged,
  input         auto_in_a_bits_user_amba_prot_secure,
  input         auto_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [3:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output        auto_out_a_bits_user_amba_prot_bufferable,
  output        auto_out_a_bits_user_amba_prot_modifiable,
  output        auto_out_a_bits_user_amba_prot_readalloc,
  output        auto_out_a_bits_user_amba_prot_writealloc,
  output        auto_out_a_bits_user_amba_prot_privileged,
  output        auto_out_a_bits_user_amba_prot_secure,
  output        auto_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum
);
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_param; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire [31:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_bufferable; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_modifiable; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_readalloc; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_writealloc; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_privileged; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_secure; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_fetch; // @[Decoupled.scala 361:21]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [31:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_bufferable; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_modifiable; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_readalloc; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_writealloc; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_privileged; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_secure; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_fetch; // @[Decoupled.scala 361:21]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [29:0] bundleOut_0_a_q_io_covSum; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire [29:0] bundleIn_0_d_q_io_covSum; // @[Decoupled.scala 361:21]
  wire [29:0] TLBuffer_2_covSum;
  wire [29:0] bundleOut_0_a_q_sum;
  wire [29:0] bundleIn_0_d_q_sum;
  Queue_4 bundleOut_0_a_q ( // @[Decoupled.scala 361:21]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_user_amba_prot_bufferable(bundleOut_0_a_q_io_enq_bits_user_amba_prot_bufferable),
    .io_enq_bits_user_amba_prot_modifiable(bundleOut_0_a_q_io_enq_bits_user_amba_prot_modifiable),
    .io_enq_bits_user_amba_prot_readalloc(bundleOut_0_a_q_io_enq_bits_user_amba_prot_readalloc),
    .io_enq_bits_user_amba_prot_writealloc(bundleOut_0_a_q_io_enq_bits_user_amba_prot_writealloc),
    .io_enq_bits_user_amba_prot_privileged(bundleOut_0_a_q_io_enq_bits_user_amba_prot_privileged),
    .io_enq_bits_user_amba_prot_secure(bundleOut_0_a_q_io_enq_bits_user_amba_prot_secure),
    .io_enq_bits_user_amba_prot_fetch(bundleOut_0_a_q_io_enq_bits_user_amba_prot_fetch),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_user_amba_prot_bufferable(bundleOut_0_a_q_io_deq_bits_user_amba_prot_bufferable),
    .io_deq_bits_user_amba_prot_modifiable(bundleOut_0_a_q_io_deq_bits_user_amba_prot_modifiable),
    .io_deq_bits_user_amba_prot_readalloc(bundleOut_0_a_q_io_deq_bits_user_amba_prot_readalloc),
    .io_deq_bits_user_amba_prot_writealloc(bundleOut_0_a_q_io_deq_bits_user_amba_prot_writealloc),
    .io_deq_bits_user_amba_prot_privileged(bundleOut_0_a_q_io_deq_bits_user_amba_prot_privileged),
    .io_deq_bits_user_amba_prot_secure(bundleOut_0_a_q_io_deq_bits_user_amba_prot_secure),
    .io_deq_bits_user_amba_prot_fetch(bundleOut_0_a_q_io_deq_bits_user_amba_prot_fetch),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_covSum(bundleOut_0_a_q_io_covSum)
  );
  Queue_5 bundleIn_0_d_q ( // @[Decoupled.scala 361:21]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt),
    .io_covSum(bundleIn_0_d_q_io_covSum)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_bufferable = bundleOut_0_a_q_io_deq_bits_user_amba_prot_bufferable; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_modifiable = bundleOut_0_a_q_io_deq_bits_user_amba_prot_modifiable; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_readalloc = bundleOut_0_a_q_io_deq_bits_user_amba_prot_readalloc; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_writealloc = bundleOut_0_a_q_io_deq_bits_user_amba_prot_writealloc; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_privileged = bundleOut_0_a_q_io_deq_bits_user_amba_prot_privileged; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_secure = bundleOut_0_a_q_io_deq_bits_user_amba_prot_secure; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_fetch = bundleOut_0_a_q_io_deq_bits_user_amba_prot_fetch; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 Decoupled.scala 365:17]
  assign bundleOut_0_a_q_clock = clock;
  assign bundleOut_0_a_q_reset = reset;
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_clock = clock;
  assign bundleIn_0_d_q_reset = reset;
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBuffer_2_covSum = 30'h0;
  assign bundleOut_0_a_q_sum = TLBuffer_2_covSum + bundleOut_0_a_q_io_covSum;
  assign bundleIn_0_d_q_sum = bundleOut_0_a_q_sum + bundleIn_0_d_q_io_covSum;
  assign io_covSum = bundleIn_0_d_q_sum;
endmodule
module TLFIFOFixer_2(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [3:0]  auto_in_a_bits_size,
  input  [3:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input         auto_in_a_bits_user_amba_prot_bufferable,
  input         auto_in_a_bits_user_amba_prot_modifiable,
  input         auto_in_a_bits_user_amba_prot_readalloc,
  input         auto_in_a_bits_user_amba_prot_writealloc,
  input         auto_in_a_bits_user_amba_prot_privileged,
  input         auto_in_a_bits_user_amba_prot_secure,
  input         auto_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [3:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [3:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output        auto_out_a_bits_user_amba_prot_bufferable,
  output        auto_out_a_bits_user_amba_prot_modifiable,
  output        auto_out_a_bits_user_amba_prot_readalloc,
  output        auto_out_a_bits_user_amba_prot_writealloc,
  output        auto_out_a_bits_user_amba_prot_privileged,
  output        auto_out_a_bits_user_amba_prot_secure,
  output        auto_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] _a_id_T_1 = {1'b0,$signed(auto_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_3 = $signed(_a_id_T_1) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  a_id = $signed(_a_id_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire  a_noDomain = ~a_id; // @[FIFOFixer.scala 55:29]
  wire  stalls_a_sel = ~auto_in_a_bits_source[3]; // @[Parameters.scala 54:32]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25]
  reg  flight_0; // @[FIFOFixer.scala 71:27]
  reg  flight_1; // @[FIFOFixer.scala 71:27]
  reg  flight_2; // @[FIFOFixer.scala 71:27]
  reg  flight_3; // @[FIFOFixer.scala 71:27]
  reg  flight_4; // @[FIFOFixer.scala 71:27]
  reg  flight_5; // @[FIFOFixer.scala 71:27]
  reg  flight_6; // @[FIFOFixer.scala 71:27]
  reg  flight_7; // @[FIFOFixer.scala 71:27]
  reg  stalls_id; // @[Reg.scala 16:16]
  wire  stalls_0 = stalls_a_sel & a_first & (flight_0 | flight_1 | flight_2 | flight_3 | flight_4 | flight_5 | flight_6
     | flight_7) & (a_noDomain | stalls_id != a_id); // @[FIFOFixer.scala 80:50]
  reg  flight_8; // @[FIFOFixer.scala 71:27]
  reg  flight_9; // @[FIFOFixer.scala 71:27]
  reg  flight_10; // @[FIFOFixer.scala 71:27]
  reg  flight_11; // @[FIFOFixer.scala 71:27]
  reg  flight_12; // @[FIFOFixer.scala 71:27]
  reg  flight_13; // @[FIFOFixer.scala 71:27]
  reg  flight_14; // @[FIFOFixer.scala 71:27]
  reg  flight_15; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_1; // @[Reg.scala 16:16]
  wire  stalls_1 = auto_in_a_bits_source[3] & a_first & (flight_8 | flight_9 | flight_10 | flight_11 | flight_12 |
    flight_13 | flight_14 | flight_15) & (a_noDomain | stalls_id_1 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stall = stalls_0 | stalls_1; // @[FIFOFixer.scala 83:49]
  wire  _bundleIn_0_a_ready_T = ~stall; // @[FIFOFixer.scala 88:50]
  wire  bundleIn_0_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  wire  _a_first_T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _a_first_beats1_decode_T_1 = 27'hfff << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [11:0] _a_first_beats1_decode_T_3 = ~_a_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] a_first_beats1_decode = _a_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28]
  wire  _d_first_T = auto_in_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28]
  wire  d_first_first = d_first_counter == 9'h0; // @[Edges.scala 230:25]
  wire  d_first = d_first_first & auto_out_d_bits_opcode != 3'h6; // @[FIFOFixer.scala 67:42]
  wire  _GEN_18 = a_first & _a_first_T ? 4'h0 == auto_in_a_bits_source | flight_0 : flight_0; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_19 = a_first & _a_first_T ? 4'h1 == auto_in_a_bits_source | flight_1 : flight_1; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_20 = a_first & _a_first_T ? 4'h2 == auto_in_a_bits_source | flight_2 : flight_2; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_21 = a_first & _a_first_T ? 4'h3 == auto_in_a_bits_source | flight_3 : flight_3; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_22 = a_first & _a_first_T ? 4'h4 == auto_in_a_bits_source | flight_4 : flight_4; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_23 = a_first & _a_first_T ? 4'h5 == auto_in_a_bits_source | flight_5 : flight_5; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_24 = a_first & _a_first_T ? 4'h6 == auto_in_a_bits_source | flight_6 : flight_6; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_25 = a_first & _a_first_T ? 4'h7 == auto_in_a_bits_source | flight_7 : flight_7; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_26 = a_first & _a_first_T ? 4'h8 == auto_in_a_bits_source | flight_8 : flight_8; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_27 = a_first & _a_first_T ? 4'h9 == auto_in_a_bits_source | flight_9 : flight_9; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_28 = a_first & _a_first_T ? 4'ha == auto_in_a_bits_source | flight_10 : flight_10; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_29 = a_first & _a_first_T ? 4'hb == auto_in_a_bits_source | flight_11 : flight_11; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_30 = a_first & _a_first_T ? 4'hc == auto_in_a_bits_source | flight_12 : flight_12; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_31 = a_first & _a_first_T ? 4'hd == auto_in_a_bits_source | flight_13 : flight_13; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_32 = a_first & _a_first_T ? 4'he == auto_in_a_bits_source | flight_14 : flight_14; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_33 = a_first & _a_first_T ? 4'hf == auto_in_a_bits_source | flight_15 : flight_15; // @[FIFOFixer.scala 71:27 72:37]
  wire  _stalls_id_T_1 = _a_first_T & stalls_a_sel; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_5 = _a_first_T & auto_in_a_bits_source[3]; // @[FIFOFixer.scala 77:49]
  reg [2:0] TLFIFOFixer_2_covState; // @[Register tracking TLFIFOFixer_2 state]
  reg  TLFIFOFixer_2_covMap [0:7]; // @[Coverage map for TLFIFOFixer_2]
  wire  TLFIFOFixer_2_covMap_read_en; // @[Coverage map for TLFIFOFixer_2]
  wire [2:0] TLFIFOFixer_2_covMap_read_addr; // @[Coverage map for TLFIFOFixer_2]
  wire  TLFIFOFixer_2_covMap_read_data; // @[Coverage map for TLFIFOFixer_2]
  wire  TLFIFOFixer_2_covMap_write_data; // @[Coverage map for TLFIFOFixer_2]
  wire [2:0] TLFIFOFixer_2_covMap_write_addr; // @[Coverage map for TLFIFOFixer_2]
  wire  TLFIFOFixer_2_covMap_write_mask; // @[Coverage map for TLFIFOFixer_2]
  wire  TLFIFOFixer_2_covMap_write_en; // @[Coverage map for TLFIFOFixer_2]
  reg [29:0] TLFIFOFixer_2_covSum; // @[Sum of coverage map]
  wire  stalls_id_shl;
  wire [2:0] stalls_id_pad;
  wire [1:0] stalls_id_1_shl;
  wire [2:0] stalls_id_1_pad;
  wire [2:0] flight_1_shl;
  wire [2:0] flight_1_pad;
  wire [2:0] flight_12_shl;
  wire [2:0] flight_12_pad;
  wire [2:0] flight_8_shl;
  wire [2:0] flight_8_pad;
  wire [2:0] flight_9_shl;
  wire [2:0] flight_9_pad;
  wire [2:0] flight_10_shl;
  wire [2:0] flight_10_pad;
  wire [2:0] flight_5_shl;
  wire [2:0] flight_5_pad;
  wire [2:0] flight_15_shl;
  wire [2:0] flight_15_pad;
  wire [2:0] flight_14_shl;
  wire [2:0] flight_14_pad;
  wire [2:0] flight_13_shl;
  wire [2:0] flight_13_pad;
  wire [2:0] flight_7_shl;
  wire [2:0] flight_7_pad;
  wire [2:0] flight_0_shl;
  wire [2:0] flight_0_pad;
  wire [2:0] flight_11_shl;
  wire [2:0] flight_11_pad;
  wire [2:0] flight_6_shl;
  wire [2:0] flight_6_pad;
  wire [2:0] flight_3_shl;
  wire [2:0] flight_3_pad;
  wire [2:0] flight_2_shl;
  wire [2:0] flight_2_pad;
  wire [2:0] flight_4_shl;
  wire [2:0] flight_4_pad;
  wire [2:0] TLFIFOFixer_2_xor7;
  wire [2:0] TLFIFOFixer_2_xor8;
  wire [2:0] TLFIFOFixer_2_xor3;
  wire [2:0] TLFIFOFixer_2_xor9;
  wire [2:0] TLFIFOFixer_2_xor22;
  wire [2:0] TLFIFOFixer_2_xor10;
  wire [2:0] TLFIFOFixer_2_xor4;
  wire [2:0] TLFIFOFixer_2_xor1;
  wire [2:0] TLFIFOFixer_2_xor11;
  wire [2:0] TLFIFOFixer_2_xor12;
  wire [2:0] TLFIFOFixer_2_xor5;
  wire [2:0] TLFIFOFixer_2_xor13;
  wire [2:0] TLFIFOFixer_2_xor30;
  wire [2:0] TLFIFOFixer_2_xor14;
  wire [2:0] TLFIFOFixer_2_xor6;
  wire [2:0] TLFIFOFixer_2_xor2;
  wire [2:0] TLFIFOFixer_2_xor0;
  assign auto_in_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  assign auto_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = auto_in_a_valid & _bundleIn_0_a_ready_T; // @[FIFOFixer.scala 87:33]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLFIFOFixer_2_covMap_read_en = 1'h1;
  assign TLFIFOFixer_2_covMap_read_addr = TLFIFOFixer_2_covState;
  assign TLFIFOFixer_2_covMap_read_data = TLFIFOFixer_2_covMap[TLFIFOFixer_2_covMap_read_addr]; // @[Coverage map for TLFIFOFixer_2]
  assign TLFIFOFixer_2_covMap_write_data = 1'h1;
  assign TLFIFOFixer_2_covMap_write_addr = TLFIFOFixer_2_covState;
  assign TLFIFOFixer_2_covMap_write_mask = 1'h1;
  assign TLFIFOFixer_2_covMap_write_en = ~metaReset;
  assign stalls_id_shl = stalls_id;
  assign stalls_id_pad = {2'h0,stalls_id_shl};
  assign stalls_id_1_shl = {stalls_id_1, 1'h0};
  assign stalls_id_1_pad = {1'h0,stalls_id_1_shl};
  assign flight_1_shl = {flight_1, 2'h0};
  assign flight_1_pad = flight_1_shl;
  assign flight_12_shl = {flight_12, 2'h0};
  assign flight_12_pad = flight_12_shl;
  assign flight_8_shl = {flight_8, 2'h0};
  assign flight_8_pad = flight_8_shl;
  assign flight_9_shl = {flight_9, 2'h0};
  assign flight_9_pad = flight_9_shl;
  assign flight_10_shl = {flight_10, 2'h0};
  assign flight_10_pad = flight_10_shl;
  assign flight_5_shl = {flight_5, 2'h0};
  assign flight_5_pad = flight_5_shl;
  assign flight_15_shl = {flight_15, 2'h0};
  assign flight_15_pad = flight_15_shl;
  assign flight_14_shl = {flight_14, 2'h0};
  assign flight_14_pad = flight_14_shl;
  assign flight_13_shl = {flight_13, 2'h0};
  assign flight_13_pad = flight_13_shl;
  assign flight_7_shl = {flight_7, 2'h0};
  assign flight_7_pad = flight_7_shl;
  assign flight_0_shl = {flight_0, 2'h0};
  assign flight_0_pad = flight_0_shl;
  assign flight_11_shl = {flight_11, 2'h0};
  assign flight_11_pad = flight_11_shl;
  assign flight_6_shl = {flight_6, 2'h0};
  assign flight_6_pad = flight_6_shl;
  assign flight_3_shl = {flight_3, 2'h0};
  assign flight_3_pad = flight_3_shl;
  assign flight_2_shl = {flight_2, 2'h0};
  assign flight_2_pad = flight_2_shl;
  assign flight_4_shl = {flight_4, 2'h0};
  assign flight_4_pad = flight_4_shl;
  assign TLFIFOFixer_2_xor7 = stalls_id_pad ^ stalls_id_1_pad;
  assign TLFIFOFixer_2_xor8 = flight_1_pad ^ flight_12_pad;
  assign TLFIFOFixer_2_xor3 = TLFIFOFixer_2_xor7 ^ TLFIFOFixer_2_xor8;
  assign TLFIFOFixer_2_xor9 = flight_8_pad ^ flight_9_pad;
  assign TLFIFOFixer_2_xor22 = flight_5_pad ^ flight_15_pad;
  assign TLFIFOFixer_2_xor10 = flight_10_pad ^ TLFIFOFixer_2_xor22;
  assign TLFIFOFixer_2_xor4 = TLFIFOFixer_2_xor9 ^ TLFIFOFixer_2_xor10;
  assign TLFIFOFixer_2_xor1 = TLFIFOFixer_2_xor3 ^ TLFIFOFixer_2_xor4;
  assign TLFIFOFixer_2_xor11 = flight_14_pad ^ flight_13_pad;
  assign TLFIFOFixer_2_xor12 = flight_7_pad ^ flight_0_pad;
  assign TLFIFOFixer_2_xor5 = TLFIFOFixer_2_xor11 ^ TLFIFOFixer_2_xor12;
  assign TLFIFOFixer_2_xor13 = flight_11_pad ^ flight_6_pad;
  assign TLFIFOFixer_2_xor30 = flight_2_pad ^ flight_4_pad;
  assign TLFIFOFixer_2_xor14 = flight_3_pad ^ TLFIFOFixer_2_xor30;
  assign TLFIFOFixer_2_xor6 = TLFIFOFixer_2_xor13 ^ TLFIFOFixer_2_xor14;
  assign TLFIFOFixer_2_xor2 = TLFIFOFixer_2_xor5 ^ TLFIFOFixer_2_xor6;
  assign TLFIFOFixer_2_xor0 = TLFIFOFixer_2_xor1 ^ TLFIFOFixer_2_xor2;
  assign io_covSum = TLFIFOFixer_2_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin
      if (a_first) begin
        if (a_first_beats1_opdata) begin
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_0 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h0 == auto_out_d_bits_source) begin
        flight_0 <= 1'h0;
      end else begin
        flight_0 <= _GEN_18;
      end
    end else begin
      flight_0 <= _GEN_18;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_1 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h1 == auto_out_d_bits_source) begin
        flight_1 <= 1'h0;
      end else begin
        flight_1 <= _GEN_19;
      end
    end else begin
      flight_1 <= _GEN_19;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_2 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h2 == auto_out_d_bits_source) begin
        flight_2 <= 1'h0;
      end else begin
        flight_2 <= _GEN_20;
      end
    end else begin
      flight_2 <= _GEN_20;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_3 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h3 == auto_out_d_bits_source) begin
        flight_3 <= 1'h0;
      end else begin
        flight_3 <= _GEN_21;
      end
    end else begin
      flight_3 <= _GEN_21;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_4 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h4 == auto_out_d_bits_source) begin
        flight_4 <= 1'h0;
      end else begin
        flight_4 <= _GEN_22;
      end
    end else begin
      flight_4 <= _GEN_22;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_5 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h5 == auto_out_d_bits_source) begin
        flight_5 <= 1'h0;
      end else begin
        flight_5 <= _GEN_23;
      end
    end else begin
      flight_5 <= _GEN_23;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_6 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h6 == auto_out_d_bits_source) begin
        flight_6 <= 1'h0;
      end else begin
        flight_6 <= _GEN_24;
      end
    end else begin
      flight_6 <= _GEN_24;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_7 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h7 == auto_out_d_bits_source) begin
        flight_7 <= 1'h0;
      end else begin
        flight_7 <= _GEN_25;
      end
    end else begin
      flight_7 <= _GEN_25;
    end
    if (_stalls_id_T_1) begin // @[Reg.scala 17:18]
      stalls_id <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_8 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h8 == auto_out_d_bits_source) begin
        flight_8 <= 1'h0;
      end else begin
        flight_8 <= _GEN_26;
      end
    end else begin
      flight_8 <= _GEN_26;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_9 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'h9 == auto_out_d_bits_source) begin
        flight_9 <= 1'h0;
      end else begin
        flight_9 <= _GEN_27;
      end
    end else begin
      flight_9 <= _GEN_27;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_10 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'ha == auto_out_d_bits_source) begin
        flight_10 <= 1'h0;
      end else begin
        flight_10 <= _GEN_28;
      end
    end else begin
      flight_10 <= _GEN_28;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_11 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'hb == auto_out_d_bits_source) begin
        flight_11 <= 1'h0;
      end else begin
        flight_11 <= _GEN_29;
      end
    end else begin
      flight_11 <= _GEN_29;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_12 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'hc == auto_out_d_bits_source) begin
        flight_12 <= 1'h0;
      end else begin
        flight_12 <= _GEN_30;
      end
    end else begin
      flight_12 <= _GEN_30;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_13 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'hd == auto_out_d_bits_source) begin
        flight_13 <= 1'h0;
      end else begin
        flight_13 <= _GEN_31;
      end
    end else begin
      flight_13 <= _GEN_31;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_14 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'he == auto_out_d_bits_source) begin
        flight_14 <= 1'h0;
      end else begin
        flight_14 <= _GEN_32;
      end
    end else begin
      flight_14 <= _GEN_32;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_15 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (4'hf == auto_out_d_bits_source) begin
        flight_15 <= 1'h0;
      end else begin
        flight_15 <= _GEN_33;
      end
    end else begin
      flight_15 <= _GEN_33;
    end
    if (_stalls_id_T_5) begin // @[Reg.scala 17:18]
      stalls_id_1 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin
      if (d_first_first) begin
        if (d_first_beats1_opdata) begin
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    TLFIFOFixer_2_covState <= TLFIFOFixer_2_xor0;
    if (TLFIFOFixer_2_covMap_write_en & TLFIFOFixer_2_covMap_write_mask) begin
      TLFIFOFixer_2_covMap[TLFIFOFixer_2_covMap_write_addr] <= TLFIFOFixer_2_covMap_write_data; // @[Coverage map for TLFIFOFixer_2]
    end
    if (!(TLFIFOFixer_2_covMap_read_data | metaReset)) begin
      TLFIFOFixer_2_covSum <= TLFIFOFixer_2_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    TLFIFOFixer_2_covMap[initvar] = 0; //_21[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  flight_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  flight_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  flight_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  flight_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  flight_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  flight_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  flight_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  flight_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  stalls_id = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  flight_8 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  flight_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  flight_10 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  flight_11 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  flight_12 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  flight_13 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  flight_14 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  flight_15 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  stalls_id_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  d_first_counter = _RAND_19[8:0];
  _RAND_20 = {1{`RANDOM}};
  TLFIFOFixer_2_covState = 0; //_20[2:0];
  _RAND_22 = {1{`RANDOM}};
  TLFIFOFixer_2_covSum = 0; //_22[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  ram_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_resp [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_last [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  reg  Queue_8_covState; // @[Register tracking Queue_8 state]
  reg  Queue_8_covMap [0:1]; // @[Coverage map for Queue_8]
  wire  Queue_8_covMap_read_en; // @[Coverage map for Queue_8]
  wire  Queue_8_covMap_read_addr; // @[Coverage map for Queue_8]
  wire  Queue_8_covMap_read_data; // @[Coverage map for Queue_8]
  wire  Queue_8_covMap_write_data; // @[Coverage map for Queue_8]
  wire  Queue_8_covMap_write_addr; // @[Coverage map for Queue_8]
  wire  Queue_8_covMap_write_mask; // @[Coverage map for Queue_8]
  wire  Queue_8_covMap_write_en; // @[Coverage map for Queue_8]
  reg [29:0] Queue_8_covSum; // @[Sum of coverage map]
  wire  maybe_full_shl;
  wire  maybe_full_pad;
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = 1'h0;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_resp = empty ? io_enq_bits_resp : ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_last = empty ? io_enq_bits_last : ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign Queue_8_covMap_read_en = 1'h1;
  assign Queue_8_covMap_read_addr = Queue_8_covState;
  assign Queue_8_covMap_read_data = Queue_8_covMap[Queue_8_covMap_read_addr]; // @[Coverage map for Queue_8]
  assign Queue_8_covMap_write_data = 1'h1;
  assign Queue_8_covMap_write_addr = Queue_8_covState;
  assign Queue_8_covMap_write_mask = 1'h1;
  assign Queue_8_covMap_write_en = ~metaReset;
  assign maybe_full_shl = maybe_full;
  assign maybe_full_pad = maybe_full_shl;
  assign io_covSum = Queue_8_covSum;
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
    Queue_8_covState <= maybe_full_pad;
    if (Queue_8_covMap_write_en & Queue_8_covMap_write_mask) begin
      Queue_8_covMap[Queue_8_covMap_write_addr] <= Queue_8_covMap_write_data; // @[Coverage map for Queue_8]
    end
    if (!(Queue_8_covMap_read_data | metaReset)) begin
      Queue_8_covSum <= Queue_8_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_3[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Queue_8_covMap[initvar] = 0; //_6[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  Queue_8_covState = 0; //_5[0:0];
  _RAND_7 = {1{`RANDOM}};
  Queue_8_covSum = 0; //_7[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_9(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [1:0]  io_enq_bits_resp,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [1:0]  io_deq_bits_resp,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  ram_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_resp [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_10 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_10 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  reg  Queue_9_covState; // @[Register tracking Queue_9 state]
  reg  Queue_9_covMap [0:1]; // @[Coverage map for Queue_9]
  wire  Queue_9_covMap_read_en; // @[Coverage map for Queue_9]
  wire  Queue_9_covMap_read_addr; // @[Coverage map for Queue_9]
  wire  Queue_9_covMap_read_data; // @[Coverage map for Queue_9]
  wire  Queue_9_covMap_write_data; // @[Coverage map for Queue_9]
  wire  Queue_9_covMap_write_addr; // @[Coverage map for Queue_9]
  wire  Queue_9_covMap_write_mask; // @[Coverage map for Queue_9]
  wire  Queue_9_covMap_write_en; // @[Coverage map for Queue_9]
  reg [29:0] Queue_9_covSum; // @[Sum of coverage map]
  wire  maybe_full_shl;
  wire  maybe_full_pad;
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = 1'h0;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_resp = empty ? io_enq_bits_resp : ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign Queue_9_covMap_read_en = 1'h1;
  assign Queue_9_covMap_read_addr = Queue_9_covState;
  assign Queue_9_covMap_read_data = Queue_9_covMap[Queue_9_covMap_read_addr]; // @[Coverage map for Queue_9]
  assign Queue_9_covMap_write_data = 1'h1;
  assign Queue_9_covMap_write_addr = Queue_9_covState;
  assign Queue_9_covMap_write_mask = 1'h1;
  assign Queue_9_covMap_write_en = ~metaReset;
  assign maybe_full_shl = maybe_full;
  assign maybe_full_pad = maybe_full_shl;
  assign io_covSum = Queue_9_covSum;
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
    Queue_9_covState <= maybe_full_pad;
    if (Queue_9_covMap_write_en & Queue_9_covMap_write_mask) begin
      Queue_9_covMap[Queue_9_covMap_write_addr] <= Queue_9_covMap_write_data; // @[Coverage map for Queue_9]
    end
    if (!(Queue_9_covMap_read_data | metaReset)) begin
      Queue_9_covSum <= Queue_9_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = _RAND_1[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Queue_9_covMap[initvar] = 0; //_4[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  Queue_9_covState = 0; //_3[0:0];
  _RAND_5 = {1{`RANDOM}};
  Queue_9_covSum = 0; //_5[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4ToTL(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [3:0]  auto_out_a_bits_size,
  output [3:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output        auto_out_a_bits_user_amba_prot_bufferable,
  output        auto_out_a_bits_user_amba_prot_modifiable,
  output        auto_out_a_bits_user_amba_prot_readalloc,
  output        auto_out_a_bits_user_amba_prot_writealloc,
  output        auto_out_a_bits_user_amba_prot_privileged,
  output        auto_out_a_bits_user_amba_prot_secure,
  output        auto_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [3:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  deq_clock; // @[Decoupled.scala 361:21]
  wire  deq_reset; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_bits_id; // @[Decoupled.scala 361:21]
  wire [63:0] deq_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire [1:0] deq_io_enq_bits_resp; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_bits_last; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [63:0] deq_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [1:0] deq_io_deq_bits_resp; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_bits_last; // @[Decoupled.scala 361:21]
  wire [29:0] deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  deq_metaReset; // @[Decoupled.scala 361:21]
  wire  q_b_deq_clock; // @[Decoupled.scala 361:21]
  wire  q_b_deq_reset; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_enq_bits_id; // @[Decoupled.scala 361:21]
  wire [1:0] q_b_deq_io_enq_bits_resp; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [1:0] q_b_deq_io_deq_bits_resp; // @[Decoupled.scala 361:21]
  wire [29:0] q_b_deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  q_b_deq_metaReset; // @[Decoupled.scala 361:21]
  wire [15:0] _r_size1_T = {auto_in_ar_bits_len,8'hff}; // @[Cat.scala 31:58]
  wire [22:0] _GEN_0 = {{7'd0}, _r_size1_T}; // @[Bundles.scala 31:21]
  wire [22:0] _r_size1_T_1 = _GEN_0 << auto_in_ar_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] r_size1 = _r_size1_T_1[22:8]; // @[Bundles.scala 31:30]
  wire [15:0] _r_size_T = {r_size1, 1'h0}; // @[package.scala 232:35]
  wire [15:0] _r_size_T_1 = _r_size_T | 16'h1; // @[package.scala 232:40]
  wire [15:0] _r_size_T_2 = {1'h0,r_size1}; // @[Cat.scala 31:58]
  wire [15:0] _r_size_T_3 = ~_r_size_T_2; // @[package.scala 232:53]
  wire [15:0] _r_size_T_4 = _r_size_T_1 & _r_size_T_3; // @[package.scala 232:51]
  wire [7:0] r_size_hi = _r_size_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] r_size_lo = _r_size_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  _r_size_T_5 = |r_size_hi; // @[OneHot.scala 32:14]
  wire [7:0] _r_size_T_6 = r_size_hi | r_size_lo; // @[OneHot.scala 32:28]
  wire [3:0] r_size_hi_1 = _r_size_T_6[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] r_size_lo_1 = _r_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _r_size_T_7 = |r_size_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _r_size_T_8 = r_size_hi_1 | r_size_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] r_size_hi_2 = _r_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] r_size_lo_2 = _r_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _r_size_T_9 = |r_size_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _r_size_T_10 = r_size_hi_2 | r_size_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] r_size = {_r_size_T_5,_r_size_T_7,_r_size_T_9,_r_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  _r_ok_T_1 = r_size <= 4'hc; // @[Parameters.scala 92:42]
  wire [31:0] _r_ok_T_4 = auto_in_ar_bits_addr ^ 32'h3000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_5 = {1'b0,$signed(_r_ok_T_4)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_7 = $signed(_r_ok_T_5) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_8 = $signed(_r_ok_T_7) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _r_ok_T_9 = _r_ok_T_1 & _r_ok_T_8; // @[Parameters.scala 670:56]
  wire  _r_ok_T_11 = r_size <= 4'h6; // @[Parameters.scala 92:42]
  wire [32:0] _r_ok_T_15 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_17 = $signed(_r_ok_T_15) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_18 = $signed(_r_ok_T_17) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_19 = auto_in_ar_bits_addr ^ 32'h10000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_20 = {1'b0,$signed(_r_ok_T_19)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_22 = $signed(_r_ok_T_20) & -33'sh10000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_23 = $signed(_r_ok_T_22) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_24 = auto_in_ar_bits_addr ^ 32'h20000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_25 = {1'b0,$signed(_r_ok_T_24)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_27 = $signed(_r_ok_T_25) & -33'sh2000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_28 = $signed(_r_ok_T_27) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_29 = auto_in_ar_bits_addr ^ 32'h2000000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_30 = {1'b0,$signed(_r_ok_T_29)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_32 = $signed(_r_ok_T_30) & -33'sh10000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_33 = $signed(_r_ok_T_32) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_34 = auto_in_ar_bits_addr ^ 32'hc000000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_35 = {1'b0,$signed(_r_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_37 = $signed(_r_ok_T_35) & -33'sh4000000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_38 = $signed(_r_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_39 = auto_in_ar_bits_addr ^ 32'h64000000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_40 = {1'b0,$signed(_r_ok_T_39)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_42 = $signed(_r_ok_T_40) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_43 = $signed(_r_ok_T_42) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_44 = auto_in_ar_bits_addr ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_45 = {1'b0,$signed(_r_ok_T_44)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_47 = $signed(_r_ok_T_45) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_48 = $signed(_r_ok_T_47) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _r_ok_T_54 = _r_ok_T_18 | _r_ok_T_23 | _r_ok_T_28 | _r_ok_T_33 | _r_ok_T_38 | _r_ok_T_43 | _r_ok_T_48; // @[Parameters.scala 671:42]
  wire  _r_ok_T_55 = _r_ok_T_11 & _r_ok_T_54; // @[Parameters.scala 670:56]
  wire  r_ok = _r_ok_T_9 | _r_ok_T_55; // @[Parameters.scala 672:30]
  wire [13:0] _GEN_16 = {{11'd0}, auto_in_ar_bits_addr[2:0]}; // @[ToTL.scala 90:59]
  wire [13:0] _r_addr_T_1 = 14'h3000 | _GEN_16; // @[ToTL.scala 90:59]
  wire [31:0] r_addr = r_ok ? auto_in_ar_bits_addr : {{18'd0}, _r_addr_T_1}; // @[ToTL.scala 90:23]
  reg [2:0] r_count_0; // @[ToTL.scala 91:28]
  reg [2:0] r_count_1; // @[ToTL.scala 91:28]
  wire [2:0] _GEN_1 = auto_in_ar_bits_id ? r_count_1 : r_count_0; // @[ToTL.scala 95:{50,50}]
  wire [3:0] r_id = {auto_in_ar_bits_id,_GEN_1[1:0],1'h0}; // @[Cat.scala 31:58]
  wire [29:0] _T_2 = 30'h7fff << r_size; // @[package.scala 234:77]
  wire [14:0] _T_4 = ~_T_2[14:0]; // @[package.scala 234:46]
  wire  _T_8 = ~reset; // @[ToTL.scala 98:14]
  wire [1:0] a_mask_sizeOH_shiftAmount = r_size[1:0]; // @[OneHot.scala 63:49]
  wire [3:0] _a_mask_sizeOH_T_1 = 4'h1 << a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [2:0] a_mask_sizeOH = _a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _a_mask_T = r_size >= 4'h3; // @[Misc.scala 205:21]
  wire  a_mask_size = a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  a_mask_bit = r_addr[2]; // @[Misc.scala 209:26]
  wire  a_mask_nbit = ~a_mask_bit; // @[Misc.scala 210:20]
  wire  a_mask_acc = _a_mask_T | a_mask_size & a_mask_nbit; // @[Misc.scala 214:29]
  wire  a_mask_acc_1 = _a_mask_T | a_mask_size & a_mask_bit; // @[Misc.scala 214:29]
  wire  a_mask_size_1 = a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  a_mask_bit_1 = r_addr[1]; // @[Misc.scala 209:26]
  wire  a_mask_nbit_1 = ~a_mask_bit_1; // @[Misc.scala 210:20]
  wire  a_mask_eq_2 = a_mask_nbit & a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_2 = a_mask_acc | a_mask_size_1 & a_mask_eq_2; // @[Misc.scala 214:29]
  wire  a_mask_eq_3 = a_mask_nbit & a_mask_bit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_3 = a_mask_acc | a_mask_size_1 & a_mask_eq_3; // @[Misc.scala 214:29]
  wire  a_mask_eq_4 = a_mask_bit & a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_4 = a_mask_acc_1 | a_mask_size_1 & a_mask_eq_4; // @[Misc.scala 214:29]
  wire  a_mask_eq_5 = a_mask_bit & a_mask_bit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_5 = a_mask_acc_1 | a_mask_size_1 & a_mask_eq_5; // @[Misc.scala 214:29]
  wire  a_mask_size_2 = a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  a_mask_bit_2 = r_addr[0]; // @[Misc.scala 209:26]
  wire  a_mask_nbit_2 = ~a_mask_bit_2; // @[Misc.scala 210:20]
  wire  a_mask_eq_6 = a_mask_eq_2 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_6 = a_mask_acc_2 | a_mask_size_2 & a_mask_eq_6; // @[Misc.scala 214:29]
  wire  a_mask_eq_7 = a_mask_eq_2 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_7 = a_mask_acc_2 | a_mask_size_2 & a_mask_eq_7; // @[Misc.scala 214:29]
  wire  a_mask_eq_8 = a_mask_eq_3 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_8 = a_mask_acc_3 | a_mask_size_2 & a_mask_eq_8; // @[Misc.scala 214:29]
  wire  a_mask_eq_9 = a_mask_eq_3 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_9 = a_mask_acc_3 | a_mask_size_2 & a_mask_eq_9; // @[Misc.scala 214:29]
  wire  a_mask_eq_10 = a_mask_eq_4 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_10 = a_mask_acc_4 | a_mask_size_2 & a_mask_eq_10; // @[Misc.scala 214:29]
  wire  a_mask_eq_11 = a_mask_eq_4 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_11 = a_mask_acc_4 | a_mask_size_2 & a_mask_eq_11; // @[Misc.scala 214:29]
  wire  a_mask_eq_12 = a_mask_eq_5 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_12 = a_mask_acc_5 | a_mask_size_2 & a_mask_eq_12; // @[Misc.scala 214:29]
  wire  a_mask_eq_13 = a_mask_eq_5 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_13 = a_mask_acc_5 | a_mask_size_2 & a_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] a_mask = {a_mask_acc_13,a_mask_acc_12,a_mask_acc_11,a_mask_acc_10,a_mask_acc_9,a_mask_acc_8,a_mask_acc_7,
    a_mask_acc_6}; // @[Cat.scala 31:58]
  wire  r_out_bits_user_amba_prot_privileged = auto_in_ar_bits_prot[0]; // @[ToTL.scala 105:45]
  wire  r_out_bits_user_amba_prot_secure = ~auto_in_ar_bits_prot[1]; // @[ToTL.scala 106:29]
  wire  r_out_bits_user_amba_prot_fetch = auto_in_ar_bits_prot[2]; // @[ToTL.scala 107:45]
  wire  r_out_bits_user_amba_prot_bufferable = auto_in_ar_bits_cache[0]; // @[ToTL.scala 108:46]
  wire  r_out_bits_user_amba_prot_modifiable = auto_in_ar_bits_cache[1]; // @[ToTL.scala 109:46]
  wire  r_out_bits_user_amba_prot_readalloc = auto_in_ar_bits_cache[2]; // @[ToTL.scala 110:46]
  wire  r_out_bits_user_amba_prot_writealloc = auto_in_ar_bits_cache[3]; // @[ToTL.scala 111:46]
  wire [1:0] r_sel = 2'h1 << auto_in_ar_bits_id; // @[OneHot.scala 64:12]
  reg [7:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 8'h0; // @[Arbiter.scala 88:28]
  wire  w_out_valid = auto_in_aw_valid & auto_in_w_valid; // @[ToTL.scala 135:34]
  wire [1:0] readys_valid = {w_out_valid,auto_in_ar_valid}; // @[Cat.scala 31:58]
  reg [1:0] readys_mask; // @[Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 24:30]
  wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter = {_readys_filter_T_1,w_out_valid,auto_in_ar_valid}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_17 = {{1'd0}, readys_filter[3:1]}; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_17; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_18 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready = _GEN_18 | _readys_unready_T_4; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 26:18]
  wire  readys_0 = readys_readys[0]; // @[Arbiter.scala 95:86]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  out_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 123:31]
  wire  _T_12 = out_ready & auto_in_ar_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _r_count_0_T_1 = r_count_0 + 3'h1; // @[ToTL.scala 116:43]
  wire [2:0] _r_count_1_T_1 = r_count_1 + 3'h1; // @[ToTL.scala 116:43]
  wire [15:0] _w_size1_T = {auto_in_aw_bits_len,8'hff}; // @[Cat.scala 31:58]
  wire [22:0] _GEN_30 = {{7'd0}, _w_size1_T}; // @[Bundles.scala 31:21]
  wire [22:0] _w_size1_T_1 = _GEN_30 << auto_in_aw_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] w_size1 = _w_size1_T_1[22:8]; // @[Bundles.scala 31:30]
  wire [15:0] _w_size_T = {w_size1, 1'h0}; // @[package.scala 232:35]
  wire [15:0] _w_size_T_1 = _w_size_T | 16'h1; // @[package.scala 232:40]
  wire [15:0] _w_size_T_2 = {1'h0,w_size1}; // @[Cat.scala 31:58]
  wire [15:0] _w_size_T_3 = ~_w_size_T_2; // @[package.scala 232:53]
  wire [15:0] _w_size_T_4 = _w_size_T_1 & _w_size_T_3; // @[package.scala 232:51]
  wire [7:0] w_size_hi = _w_size_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] w_size_lo = _w_size_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  _w_size_T_5 = |w_size_hi; // @[OneHot.scala 32:14]
  wire [7:0] _w_size_T_6 = w_size_hi | w_size_lo; // @[OneHot.scala 32:28]
  wire [3:0] w_size_hi_1 = _w_size_T_6[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] w_size_lo_1 = _w_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _w_size_T_7 = |w_size_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _w_size_T_8 = w_size_hi_1 | w_size_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] w_size_hi_2 = _w_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] w_size_lo_2 = _w_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _w_size_T_9 = |w_size_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _w_size_T_10 = w_size_hi_2 | w_size_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] w_size = {_w_size_T_5,_w_size_T_7,_w_size_T_9,_w_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  _w_ok_T_1 = w_size <= 4'hc; // @[Parameters.scala 92:42]
  wire [31:0] _w_ok_T_4 = auto_in_aw_bits_addr ^ 32'h3000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_5 = {1'b0,$signed(_w_ok_T_4)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_7 = $signed(_w_ok_T_5) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_8 = $signed(_w_ok_T_7) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _w_ok_T_9 = _w_ok_T_1 & _w_ok_T_8; // @[Parameters.scala 670:56]
  wire  _w_ok_T_11 = w_size <= 4'h6; // @[Parameters.scala 92:42]
  wire [32:0] _w_ok_T_15 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_17 = $signed(_w_ok_T_15) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_18 = $signed(_w_ok_T_17) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _w_ok_T_19 = auto_in_aw_bits_addr ^ 32'h2000000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_20 = {1'b0,$signed(_w_ok_T_19)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_22 = $signed(_w_ok_T_20) & -33'sh10000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_23 = $signed(_w_ok_T_22) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _w_ok_T_24 = auto_in_aw_bits_addr ^ 32'hc000000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_25 = {1'b0,$signed(_w_ok_T_24)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_27 = $signed(_w_ok_T_25) & -33'sh4000000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_28 = $signed(_w_ok_T_27) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _w_ok_T_29 = auto_in_aw_bits_addr ^ 32'h64000000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_30 = {1'b0,$signed(_w_ok_T_29)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_32 = $signed(_w_ok_T_30) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_33 = $signed(_w_ok_T_32) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _w_ok_T_34 = auto_in_aw_bits_addr ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_35 = {1'b0,$signed(_w_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_37 = $signed(_w_ok_T_35) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_38 = $signed(_w_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _w_ok_T_42 = _w_ok_T_18 | _w_ok_T_23 | _w_ok_T_28 | _w_ok_T_33 | _w_ok_T_38; // @[Parameters.scala 671:42]
  wire  _w_ok_T_43 = _w_ok_T_11 & _w_ok_T_42; // @[Parameters.scala 670:56]
  wire  w_ok = _w_ok_T_9 | _w_ok_T_43; // @[Parameters.scala 672:30]
  wire [13:0] _GEN_19 = {{11'd0}, auto_in_aw_bits_addr[2:0]}; // @[ToTL.scala 123:59]
  wire [13:0] _w_addr_T_1 = 14'h3000 | _GEN_19; // @[ToTL.scala 123:59]
  wire [31:0] w_addr = w_ok ? auto_in_aw_bits_addr : {{18'd0}, _w_addr_T_1}; // @[ToTL.scala 123:23]
  reg [2:0] w_count_0; // @[ToTL.scala 124:28]
  reg [2:0] w_count_1; // @[ToTL.scala 124:28]
  wire [2:0] _GEN_5 = auto_in_aw_bits_id ? w_count_1 : w_count_0; // @[ToTL.scala 128:{50,50}]
  wire [3:0] w_id = {auto_in_aw_bits_id,_GEN_5[1:0],1'h1}; // @[Cat.scala 31:58]
  wire  _T_16 = ~auto_in_aw_valid; // @[ToTL.scala 131:15]
  wire [29:0] _T_18 = 30'h7fff << w_size; // @[package.scala 234:77]
  wire [14:0] _T_20 = ~_T_18[14:0]; // @[package.scala 234:46]
  wire  readys_1 = readys_readys[1]; // @[Arbiter.scala 95:86]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 123:31]
  wire  bundleIn_0_aw_ready = out_1_ready & auto_in_w_valid & auto_in_w_bits_last; // @[ToTL.scala 133:48]
  wire  w_out_bits_user_amba_prot_privileged = auto_in_aw_bits_prot[0]; // @[ToTL.scala 141:45]
  wire  w_out_bits_user_amba_prot_secure = ~auto_in_aw_bits_prot[1]; // @[ToTL.scala 142:29]
  wire  w_out_bits_user_amba_prot_fetch = auto_in_aw_bits_prot[2]; // @[ToTL.scala 143:45]
  wire  w_out_bits_user_amba_prot_bufferable = auto_in_aw_bits_cache[0]; // @[ToTL.scala 144:46]
  wire  w_out_bits_user_amba_prot_modifiable = auto_in_aw_bits_cache[1]; // @[ToTL.scala 145:46]
  wire  w_out_bits_user_amba_prot_readalloc = auto_in_aw_bits_cache[2]; // @[ToTL.scala 146:46]
  wire  w_out_bits_user_amba_prot_writealloc = auto_in_aw_bits_cache[3]; // @[ToTL.scala 147:46]
  wire [1:0] w_sel = 2'h1 << auto_in_aw_bits_id; // @[OneHot.scala 64:12]
  wire  _T_36 = bundleIn_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _w_count_0_T_1 = w_count_0 + 3'h1; // @[ToTL.scala 152:43]
  wire [2:0] _w_count_1_T_1 = w_count_1 + 3'h1; // @[ToTL.scala 152:43]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 89:24]
  wire [1:0] _readys_mask_T = readys_readys & readys_valid; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[package.scala 244:43]
  wire  earlyWinner_0 = readys_0 & auto_in_ar_valid; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1 = readys_1 & w_out_valid; // @[Arbiter.scala 97:79]
  wire  _T_50 = auto_in_ar_valid | w_out_valid; // @[Arbiter.scala 107:36]
  wire  _T_51 = ~(auto_in_ar_valid | w_out_valid); // @[Arbiter.scala 107:15]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & auto_in_ar_valid | state_1 & w_out_valid; // @[Mux.scala 27:73]
  wire  sink_ACancel_earlyValid = idle ? _T_50 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [7:0] _GEN_20 = {{7'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [7:0] _beatsLeft_T_4 = beatsLeft - _GEN_20; // @[Arbiter.scala 113:52]
  wire [7:0] _T_70 = muxStateEarly_0 ? a_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_71 = muxStateEarly_1 ? auto_in_w_bits_strb : 8'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_94 = muxStateEarly_0 ? r_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_95 = muxStateEarly_1 ? w_addr : 32'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_97 = muxStateEarly_0 ? r_id : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_98 = muxStateEarly_1 ? w_id : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_100 = muxStateEarly_0 ? r_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_101 = muxStateEarly_1 ? w_size : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_106 = muxStateEarly_0 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_107 = muxStateEarly_1 ? 3'h1 : 3'h0; // @[Mux.scala 27:73]
  wire  d_hasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  ok_r_ready = deq_io_enq_ready; // @[ToTL.scala 158:23 Decoupled.scala 365:17]
  wire  ok_b_ready = q_b_deq_io_enq_ready; // @[ToTL.scala 157:23 Decoupled.scala 365:17]
  wire  bundleOut_0_d_ready = d_hasData ? ok_r_ready : ok_b_ready; // @[ToTL.scala 164:25]
  wire  _d_last_T = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _d_last_beats1_decode_T_1 = 27'hfff << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [11:0] _d_last_beats1_decode_T_3 = ~_d_last_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] d_last_beats1_decode = _d_last_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire [8:0] d_last_beats1 = d_hasData ? d_last_beats1_decode : 9'h0; // @[Edges.scala 220:14]
  reg [8:0] d_last_counter; // @[Edges.scala 228:27]
  wire [8:0] d_last_counter1 = d_last_counter - 9'h1; // @[Edges.scala 229:28]
  wire  d_last_first = d_last_counter == 9'h0; // @[Edges.scala 230:25]
  reg [2:0] b_count_0; // @[ToTL.scala 186:28]
  reg [2:0] b_count_1; // @[ToTL.scala 186:28]
  wire  q_b_bits_id = q_b_deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  wire [2:0] _GEN_11 = q_b_bits_id ? b_count_1 : b_count_0; // @[ToTL.scala 187:{43,43}]
  wire [2:0] _GEN_13 = q_b_bits_id ? w_count_1 : w_count_0; // @[ToTL.scala 187:{43,43}]
  wire  b_allow = _GEN_11 != _GEN_13; // @[ToTL.scala 187:43]
  wire [1:0] b_sel = 2'h1 << q_b_bits_id; // @[OneHot.scala 64:12]
  wire  q_b_valid = q_b_deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  wire  bundleIn_0_b_valid = q_b_valid & b_allow; // @[ToTL.scala 195:31]
  wire  _T_111 = auto_in_b_ready & bundleIn_0_b_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _b_count_0_T_1 = b_count_0 + 3'h1; // @[ToTL.scala 191:42]
  wire [2:0] _b_count_1_T_1 = b_count_1 + 3'h1; // @[ToTL.scala 191:42]
  reg [8:0] AXI4ToTL_covState; // @[Register tracking AXI4ToTL state]
  reg  AXI4ToTL_covMap [0:511]; // @[Coverage map for AXI4ToTL]
  wire  AXI4ToTL_covMap_read_en; // @[Coverage map for AXI4ToTL]
  wire [8:0] AXI4ToTL_covMap_read_addr; // @[Coverage map for AXI4ToTL]
  wire  AXI4ToTL_covMap_read_data; // @[Coverage map for AXI4ToTL]
  wire  AXI4ToTL_covMap_write_data; // @[Coverage map for AXI4ToTL]
  wire [8:0] AXI4ToTL_covMap_write_addr; // @[Coverage map for AXI4ToTL]
  wire  AXI4ToTL_covMap_write_mask; // @[Coverage map for AXI4ToTL]
  wire  AXI4ToTL_covMap_write_en; // @[Coverage map for AXI4ToTL]
  reg [29:0] AXI4ToTL_covSum; // @[Sum of coverage map]
  wire [1:0] readys_mask_shl;
  wire [8:0] readys_mask_pad;
  wire [8:0] b_count_0_shl;
  wire [8:0] b_count_0_pad;
  wire [4:0] w_count_1_shl;
  wire [8:0] w_count_1_pad;
  wire [5:0] state_1_shl;
  wire [8:0] state_1_pad;
  wire [5:0] state_0_shl;
  wire [8:0] state_0_pad;
  wire [4:0] w_count_0_shl;
  wire [8:0] w_count_0_pad;
  wire [8:0] b_count_1_shl;
  wire [8:0] b_count_1_pad;
  wire [8:0] AXI4ToTL_xor4;
  wire [8:0] AXI4ToTL_xor1;
  wire [8:0] AXI4ToTL_xor5;
  wire [8:0] AXI4ToTL_xor6;
  wire [8:0] AXI4ToTL_xor2;
  wire [8:0] AXI4ToTL_xor0;
  wire [29:0] deq_sum;
  wire [29:0] q_b_deq_sum;
  Queue_8 deq ( // @[Decoupled.scala 361:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_id(deq_io_enq_bits_id),
    .io_enq_bits_data(deq_io_enq_bits_data),
    .io_enq_bits_resp(deq_io_enq_bits_resp),
    .io_enq_bits_last(deq_io_enq_bits_last),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_id(deq_io_deq_bits_id),
    .io_deq_bits_data(deq_io_deq_bits_data),
    .io_deq_bits_resp(deq_io_deq_bits_resp),
    .io_deq_bits_last(deq_io_deq_bits_last),
    .io_covSum(deq_io_covSum),
    .metaReset(deq_metaReset)
  );
  Queue_9 q_b_deq ( // @[Decoupled.scala 361:21]
    .clock(q_b_deq_clock),
    .reset(q_b_deq_reset),
    .io_enq_ready(q_b_deq_io_enq_ready),
    .io_enq_valid(q_b_deq_io_enq_valid),
    .io_enq_bits_id(q_b_deq_io_enq_bits_id),
    .io_enq_bits_resp(q_b_deq_io_enq_bits_resp),
    .io_deq_ready(q_b_deq_io_deq_ready),
    .io_deq_valid(q_b_deq_io_deq_valid),
    .io_deq_bits_id(q_b_deq_io_deq_bits_id),
    .io_deq_bits_resp(q_b_deq_io_deq_bits_resp),
    .io_covSum(q_b_deq_io_covSum),
    .metaReset(q_b_deq_metaReset)
  );
  assign auto_in_aw_ready = out_1_ready & auto_in_w_valid & auto_in_w_bits_last; // @[ToTL.scala 133:48]
  assign auto_in_w_ready = out_1_ready & auto_in_aw_valid; // @[ToTL.scala 134:34]
  assign auto_in_b_valid = q_b_valid & b_allow; // @[ToTL.scala 195:31]
  assign auto_in_b_bits_id = q_b_deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_b_bits_resp = q_b_deq_io_deq_bits_resp; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_ar_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 123:31]
  assign auto_in_r_valid = deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  assign auto_in_r_bits_id = deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_r_bits_data = deq_io_deq_bits_data; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_r_bits_resp = deq_io_deq_bits_resp; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_r_bits_last = deq_io_deq_bits_last; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_a_valid = idle ? _T_50 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_out_a_bits_opcode = _T_106 | _T_107; // @[Mux.scala 27:73]
  assign auto_out_a_bits_size = _T_100 | _T_101; // @[Mux.scala 27:73]
  assign auto_out_a_bits_source = _T_97 | _T_98; // @[Mux.scala 27:73]
  assign auto_out_a_bits_address = _T_94 | _T_95; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_bufferable = muxStateEarly_0 & r_out_bits_user_amba_prot_bufferable |
    muxStateEarly_1 & w_out_bits_user_amba_prot_bufferable; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_modifiable = muxStateEarly_0 & r_out_bits_user_amba_prot_modifiable |
    muxStateEarly_1 & w_out_bits_user_amba_prot_modifiable; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_readalloc = muxStateEarly_0 & r_out_bits_user_amba_prot_readalloc |
    muxStateEarly_1 & w_out_bits_user_amba_prot_readalloc; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_writealloc = muxStateEarly_0 & r_out_bits_user_amba_prot_writealloc |
    muxStateEarly_1 & w_out_bits_user_amba_prot_writealloc; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_privileged = muxStateEarly_0 & r_out_bits_user_amba_prot_privileged |
    muxStateEarly_1 & w_out_bits_user_amba_prot_privileged; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_secure = muxStateEarly_0 & r_out_bits_user_amba_prot_secure | muxStateEarly_1 &
    w_out_bits_user_amba_prot_secure; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_fetch = muxStateEarly_0 & r_out_bits_user_amba_prot_fetch | muxStateEarly_1 &
    w_out_bits_user_amba_prot_fetch; // @[Mux.scala 27:73]
  assign auto_out_a_bits_mask = _T_70 | _T_71; // @[Mux.scala 27:73]
  assign auto_out_a_bits_data = muxStateEarly_1 ? auto_in_w_bits_data : 64'h0; // @[Mux.scala 27:73]
  assign auto_out_d_ready = d_hasData ? ok_r_ready : ok_b_ready; // @[ToTL.scala 164:25]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = auto_out_d_valid & d_hasData; // @[ToTL.scala 165:33]
  assign deq_io_enq_bits_id = auto_out_d_bits_source[3]; // @[ToTL.scala 168:43]
  assign deq_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign deq_io_enq_bits_resp = auto_out_d_bits_denied | auto_out_d_bits_corrupt ? 2'h2 : 2'h0; // @[ToTL.scala 160:23]
  assign deq_io_enq_bits_last = d_last_counter == 9'h1 | d_last_beats1 == 9'h0; // @[Edges.scala 231:37]
  assign deq_io_deq_ready = auto_in_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign q_b_deq_clock = clock;
  assign q_b_deq_reset = reset;
  assign q_b_deq_io_enq_valid = auto_out_d_valid & ~d_hasData; // @[ToTL.scala 166:33]
  assign q_b_deq_io_enq_bits_id = auto_out_d_bits_source[3]; // @[ToTL.scala 177:43]
  assign q_b_deq_io_enq_bits_resp = auto_out_d_bits_denied | auto_out_d_bits_corrupt ? 2'h2 : 2'h0; // @[ToTL.scala 160:23]
  assign q_b_deq_io_deq_ready = auto_in_b_ready & b_allow; // @[ToTL.scala 196:31]
  assign AXI4ToTL_covMap_read_en = 1'h1;
  assign AXI4ToTL_covMap_read_addr = AXI4ToTL_covState;
  assign AXI4ToTL_covMap_read_data = AXI4ToTL_covMap[AXI4ToTL_covMap_read_addr]; // @[Coverage map for AXI4ToTL]
  assign AXI4ToTL_covMap_write_data = 1'h1;
  assign AXI4ToTL_covMap_write_addr = AXI4ToTL_covState;
  assign AXI4ToTL_covMap_write_mask = 1'h1;
  assign AXI4ToTL_covMap_write_en = ~metaReset;
  assign readys_mask_shl = readys_mask;
  assign readys_mask_pad = {7'h0,readys_mask_shl};
  assign b_count_0_shl = {b_count_0, 6'h0};
  assign b_count_0_pad = b_count_0_shl;
  assign w_count_1_shl = {w_count_1, 2'h0};
  assign w_count_1_pad = {4'h0,w_count_1_shl};
  assign state_1_shl = {state_1, 5'h0};
  assign state_1_pad = {3'h0,state_1_shl};
  assign state_0_shl = {state_0, 5'h0};
  assign state_0_pad = {3'h0,state_0_shl};
  assign w_count_0_shl = {w_count_0, 2'h0};
  assign w_count_0_pad = {4'h0,w_count_0_shl};
  assign b_count_1_shl = {b_count_1, 6'h0};
  assign b_count_1_pad = b_count_1_shl;
  assign AXI4ToTL_xor4 = b_count_0_pad ^ w_count_1_pad;
  assign AXI4ToTL_xor1 = readys_mask_pad ^ AXI4ToTL_xor4;
  assign AXI4ToTL_xor5 = state_1_pad ^ state_0_pad;
  assign AXI4ToTL_xor6 = w_count_0_pad ^ b_count_1_pad;
  assign AXI4ToTL_xor2 = AXI4ToTL_xor5 ^ AXI4ToTL_xor6;
  assign AXI4ToTL_xor0 = AXI4ToTL_xor1 ^ AXI4ToTL_xor2;
  assign deq_sum = AXI4ToTL_covSum + deq_io_covSum;
  assign q_b_deq_sum = deq_sum + q_b_deq_io_covSum;
  assign io_covSum = q_b_deq_sum;
  assign deq_metaReset = metaReset;
  assign q_b_deq_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_0 <= 3'h0; // @[ToTL.scala 91:28]
    end else if (_T_12 & r_sel[0]) begin
      r_count_0 <= _r_count_0_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_1 <= 3'h0; // @[ToTL.scala 91:28]
    end else if (_T_12 & r_sel[1]) begin
      r_count_1 <= _r_count_1_T_1;
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 8'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin
      if (earlyWinner_1) begin
        beatsLeft <= auto_in_aw_bits_len;
      end else begin
        beatsLeft <= 8'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (latch & |readys_valid) begin
      readys_mask <= _readys_mask_T_3;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_0 <= 3'h0; // @[ToTL.scala 124:28]
    end else if (_T_36 & w_sel[0]) begin
      w_count_0 <= _w_count_0_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_1 <= 3'h0; // @[ToTL.scala 124:28]
    end else if (_T_36 & w_sel[1]) begin
      w_count_1 <= _w_count_1_T_1;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_last_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_d_last_T) begin
      if (d_last_first) begin
        if (d_hasData) begin
          d_last_counter <= d_last_beats1_decode;
        end else begin
          d_last_counter <= 9'h0;
        end
      end else begin
        d_last_counter <= d_last_counter1;
      end
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_0 <= 3'h0; // @[ToTL.scala 186:28]
    end else if (_T_111 & b_sel[0]) begin
      b_count_0 <= _b_count_0_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_1 <= 3'h0; // @[ToTL.scala 186:28]
    end else if (_T_111 & b_sel[1]) begin
      b_count_1 <= _b_count_1_T_1;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_in_ar_valid | r_size1 == _T_4) & ~reset) begin
          $fatal; // @[ToTL.scala 98:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_in_ar_valid | r_size1 == _T_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:98 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n"
            ); // @[ToTL.scala 98:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_in_aw_valid | w_size1 == _T_20) & _T_8) begin
          $fatal; // @[ToTL.scala 131:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~auto_in_aw_valid | w_size1 == _T_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:131 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n"
            ); // @[ToTL.scala 131:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_16 | auto_in_aw_bits_len == 8'h0 | auto_in_aw_bits_size == 3'h3) & _T_8) begin
          $fatal; // @[ToTL.scala 132:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(_T_16 | auto_in_aw_bits_len == 8'h0 | auto_in_aw_bits_size == 3'h3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:132 assert (!in.aw.valid || in.aw.bits.len === UInt(0) || in.aw.bits.size === UInt(log2Ceil(beatBytes))) // because aligned\n"
            ); // @[ToTL.scala 132:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & _T_8) begin
          $fatal; // @[Arbiter.scala 22:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1) & _T_8) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~earlyWinner_0 | ~earlyWinner_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(auto_in_ar_valid | w_out_valid) | (earlyWinner_0 | earlyWinner_1)) & _T_8) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~(auto_in_ar_valid | w_out_valid) | (earlyWinner_0 | earlyWinner_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_51 | _T_50) & _T_8) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(_T_51 | _T_50)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    AXI4ToTL_covState <= AXI4ToTL_xor0;
    if (AXI4ToTL_covMap_write_en & AXI4ToTL_covMap_write_mask) begin
      AXI4ToTL_covMap[AXI4ToTL_covMap_write_addr] <= AXI4ToTL_covMap_write_data; // @[Coverage map for AXI4ToTL]
    end
    if (!(AXI4ToTL_covMap_read_data | metaReset)) begin
      AXI4ToTL_covSum <= AXI4ToTL_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    AXI4ToTL_covMap[initvar] = 0; //_12[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_count_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  r_count_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  beatsLeft = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  readys_mask = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  state_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  w_count_0 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  w_count_1 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  state_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  d_last_counter = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  b_count_0 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  b_count_1 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  AXI4ToTL_covState = 0; //_11[8:0];
  _RAND_13 = {1{`RANDOM}};
  AXI4ToTL_covSum = 0; //_13[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QueueCompatibility(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [6:0]  io_enq_bits_extra_id,
  input         io_enq_bits_real_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [6:0]  io_deq_bits_extra_id,
  output        io_deq_bits_real_last,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [6:0] ram_extra_id [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [6:0] ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [6:0] ram_extra_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_extra_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_extra_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_extra_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_real_last [0:3]; // @[Decoupled.scala 259:95]
  wire  ram_real_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_real_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_real_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_real_last_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_real_last_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_real_last_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_real_last_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  wire [29:0] QueueCompatibility_covSum;
  assign ram_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_extra_id_MPORT_data = io_enq_bits_extra_id;
  assign ram_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_extra_id_MPORT_mask = 1'h1;
  assign ram_extra_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_real_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_real_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_real_last_io_deq_bits_MPORT_data = ram_real_last[ram_real_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_real_last_MPORT_data = io_enq_bits_real_last;
  assign ram_real_last_MPORT_addr = enq_ptr_value;
  assign ram_real_last_MPORT_mask = 1'h1;
  assign ram_real_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_extra_id = ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_real_last = ram_real_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign QueueCompatibility_covSum = 30'h0;
  assign io_covSum = QueueCompatibility_covSum;
  always @(posedge clock) begin
    if (ram_extra_id_MPORT_en & ram_extra_id_MPORT_mask) begin
      ram_extra_id[ram_extra_id_MPORT_addr] <= ram_extra_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_real_last_MPORT_en & ram_real_last_MPORT_mask) begin
      ram_real_last[ram_real_last_MPORT_addr] <= ram_real_last_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      enq_ptr_value <= _value_T_1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      deq_ptr_value <= _value_T_3;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_extra_id[initvar] = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_real_last[initvar] = _RAND_1[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4UserYanker(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [6:0]  auto_in_aw_bits_echo_extra_id,
  input         auto_in_aw_bits_echo_real_last,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [6:0]  auto_in_b_bits_echo_extra_id,
  output        auto_in_b_bits_echo_real_last,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [6:0]  auto_in_ar_bits_echo_extra_id,
  input         auto_in_ar_bits_echo_real_last,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [6:0]  auto_in_r_bits_echo_extra_id,
  output        auto_in_r_bits_echo_real_last,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last,
  output [29:0] io_covSum
);
  wire  QueueCompatibility_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_1_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_1_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_1_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_2_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_2_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_2_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_3_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [6:0] QueueCompatibility_3_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_3_io_covSum; // @[UserYanker.scala 47:17]
  wire  _ar_ready_WIRE_0 = QueueCompatibility_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _ar_ready_WIRE_1 = QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_1 = auto_in_ar_bits_id ? _ar_ready_WIRE_1 : _ar_ready_WIRE_0; // @[UserYanker.scala 56:{36,36}]
  wire  _r_valid_WIRE_0 = QueueCompatibility_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _r_valid_WIRE_1 = QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_3 = auto_out_r_bits_id ? _r_valid_WIRE_1 : _r_valid_WIRE_0; // @[UserYanker.scala 63:{28,28}]
  wire  _T_3 = ~reset; // @[UserYanker.scala 63:14]
  wire  _r_bits_WIRE_0_real_last = QueueCompatibility_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _r_bits_WIRE_1_real_last = QueueCompatibility_1_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire [6:0] _r_bits_WIRE_0_extra_id = QueueCompatibility_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [6:0] _r_bits_WIRE_1_extra_id = QueueCompatibility_1_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [1:0] _arsel_T = 2'h1 << auto_in_ar_bits_id; // @[OneHot.scala 64:12]
  wire  arsel_0 = _arsel_T[0]; // @[UserYanker.scala 67:55]
  wire  arsel_1 = _arsel_T[1]; // @[UserYanker.scala 67:55]
  wire [1:0] _rsel_T = 2'h1 << auto_out_r_bits_id; // @[OneHot.scala 64:12]
  wire  rsel_0 = _rsel_T[0]; // @[UserYanker.scala 68:55]
  wire  rsel_1 = _rsel_T[1]; // @[UserYanker.scala 68:55]
  wire  _aw_ready_WIRE_0 = QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _aw_ready_WIRE_1 = QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_9 = auto_in_aw_bits_id ? _aw_ready_WIRE_1 : _aw_ready_WIRE_0; // @[UserYanker.scala 77:{36,36}]
  wire  _b_valid_WIRE_0 = QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _b_valid_WIRE_1 = QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_11 = auto_out_b_bits_id ? _b_valid_WIRE_1 : _b_valid_WIRE_0; // @[UserYanker.scala 84:{28,28}]
  wire  _b_bits_WIRE_0_real_last = QueueCompatibility_2_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _b_bits_WIRE_1_real_last = QueueCompatibility_3_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire [6:0] _b_bits_WIRE_0_extra_id = QueueCompatibility_2_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [6:0] _b_bits_WIRE_1_extra_id = QueueCompatibility_3_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [1:0] _awsel_T = 2'h1 << auto_in_aw_bits_id; // @[OneHot.scala 64:12]
  wire  awsel_0 = _awsel_T[0]; // @[UserYanker.scala 88:55]
  wire  awsel_1 = _awsel_T[1]; // @[UserYanker.scala 88:55]
  wire [1:0] _bsel_T = 2'h1 << auto_out_b_bits_id; // @[OneHot.scala 64:12]
  wire  bsel_0 = _bsel_T[0]; // @[UserYanker.scala 89:55]
  wire  bsel_1 = _bsel_T[1]; // @[UserYanker.scala 89:55]
  wire [29:0] AXI4UserYanker_covSum;
  wire [29:0] QueueCompatibility_sum;
  wire [29:0] QueueCompatibility_1_sum;
  wire [29:0] QueueCompatibility_2_sum;
  wire [29:0] QueueCompatibility_3_sum;
  QueueCompatibility QueueCompatibility ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_clock),
    .reset(QueueCompatibility_reset),
    .io_enq_ready(QueueCompatibility_io_enq_ready),
    .io_enq_valid(QueueCompatibility_io_enq_valid),
    .io_enq_bits_extra_id(QueueCompatibility_io_enq_bits_extra_id),
    .io_enq_bits_real_last(QueueCompatibility_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_io_deq_ready),
    .io_deq_valid(QueueCompatibility_io_deq_valid),
    .io_deq_bits_extra_id(QueueCompatibility_io_deq_bits_extra_id),
    .io_deq_bits_real_last(QueueCompatibility_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_io_covSum)
  );
  QueueCompatibility QueueCompatibility_1 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_1_clock),
    .reset(QueueCompatibility_1_reset),
    .io_enq_ready(QueueCompatibility_1_io_enq_ready),
    .io_enq_valid(QueueCompatibility_1_io_enq_valid),
    .io_enq_bits_extra_id(QueueCompatibility_1_io_enq_bits_extra_id),
    .io_enq_bits_real_last(QueueCompatibility_1_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_1_io_deq_ready),
    .io_deq_valid(QueueCompatibility_1_io_deq_valid),
    .io_deq_bits_extra_id(QueueCompatibility_1_io_deq_bits_extra_id),
    .io_deq_bits_real_last(QueueCompatibility_1_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_1_io_covSum)
  );
  QueueCompatibility QueueCompatibility_2 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_2_clock),
    .reset(QueueCompatibility_2_reset),
    .io_enq_ready(QueueCompatibility_2_io_enq_ready),
    .io_enq_valid(QueueCompatibility_2_io_enq_valid),
    .io_enq_bits_extra_id(QueueCompatibility_2_io_enq_bits_extra_id),
    .io_enq_bits_real_last(QueueCompatibility_2_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_2_io_deq_ready),
    .io_deq_valid(QueueCompatibility_2_io_deq_valid),
    .io_deq_bits_extra_id(QueueCompatibility_2_io_deq_bits_extra_id),
    .io_deq_bits_real_last(QueueCompatibility_2_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_2_io_covSum)
  );
  QueueCompatibility QueueCompatibility_3 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_3_clock),
    .reset(QueueCompatibility_3_reset),
    .io_enq_ready(QueueCompatibility_3_io_enq_ready),
    .io_enq_valid(QueueCompatibility_3_io_enq_valid),
    .io_enq_bits_extra_id(QueueCompatibility_3_io_enq_bits_extra_id),
    .io_enq_bits_real_last(QueueCompatibility_3_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_3_io_deq_ready),
    .io_deq_valid(QueueCompatibility_3_io_deq_valid),
    .io_deq_bits_extra_id(QueueCompatibility_3_io_deq_bits_extra_id),
    .io_deq_bits_real_last(QueueCompatibility_3_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_3_io_covSum)
  );
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_9; // @[UserYanker.scala 77:36]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_echo_extra_id = auto_out_b_bits_id ? _b_bits_WIRE_1_extra_id : _b_bits_WIRE_0_extra_id; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_b_bits_echo_real_last = auto_out_b_bits_id ? _b_bits_WIRE_1_real_last : _b_bits_WIRE_0_real_last; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_1; // @[UserYanker.scala 56:36]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_echo_extra_id = auto_out_r_bits_id ? _r_bits_WIRE_1_extra_id : _r_bits_WIRE_0_extra_id; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_echo_real_last = auto_out_r_bits_id ? _r_bits_WIRE_1_real_last : _r_bits_WIRE_0_real_last; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_9; // @[UserYanker.scala 78:36]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_valid = auto_in_w_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_1; // @[UserYanker.scala 57:36]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_clock = clock;
  assign QueueCompatibility_reset = reset;
  assign QueueCompatibility_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_0; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_0 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_1_clock = clock;
  assign QueueCompatibility_1_reset = reset;
  assign QueueCompatibility_1_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_1; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_1_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_1 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_2_clock = clock;
  assign QueueCompatibility_2_reset = reset;
  assign QueueCompatibility_2_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_0; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_2_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_0; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_3_clock = clock;
  assign QueueCompatibility_3_reset = reset;
  assign QueueCompatibility_3_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_1; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_3_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_1; // @[UserYanker.scala 91:53]
  assign AXI4UserYanker_covSum = 30'h0;
  assign QueueCompatibility_sum = AXI4UserYanker_covSum + QueueCompatibility_io_covSum;
  assign QueueCompatibility_1_sum = QueueCompatibility_sum + QueueCompatibility_1_io_covSum;
  assign QueueCompatibility_2_sum = QueueCompatibility_1_sum + QueueCompatibility_2_io_covSum;
  assign QueueCompatibility_3_sum = QueueCompatibility_2_sum + QueueCompatibility_3_io_covSum;
  assign io_covSum = QueueCompatibility_3_sum;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_r_valid | _GEN_3) & ~reset) begin
          $fatal; // @[UserYanker.scala 63:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_out_r_valid | _GEN_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:63 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 63:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_b_valid | _GEN_11) & _T_3) begin
          $fatal; // @[UserYanker.scala 84:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~auto_out_b_valid | _GEN_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:84 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 84:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_10(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input  [3:0]  io_enq_bits_cache,
  input  [2:0]  io_enq_bits_prot,
  input  [6:0]  io_enq_bits_echo_extra_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [6:0]  io_deq_bits_echo_extra_id,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg  ram_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_len [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_burst [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_cache [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_cache_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_cache_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_cache_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_prot [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_prot_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_prot_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_prot_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_en; // @[Decoupled.scala 259:95]
  reg [6:0] ram_echo_extra_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_echo_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [6:0] ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [6:0] ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_echo_extra_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_echo_extra_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_echo_extra_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_18 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_18 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  reg  Queue_10_covState; // @[Register tracking Queue_10 state]
  reg  Queue_10_covMap [0:1]; // @[Coverage map for Queue_10]
  wire  Queue_10_covMap_read_en; // @[Coverage map for Queue_10]
  wire  Queue_10_covMap_read_addr; // @[Coverage map for Queue_10]
  wire  Queue_10_covMap_read_data; // @[Coverage map for Queue_10]
  wire  Queue_10_covMap_write_data; // @[Coverage map for Queue_10]
  wire  Queue_10_covMap_write_addr; // @[Coverage map for Queue_10]
  wire  Queue_10_covMap_write_mask; // @[Coverage map for Queue_10]
  wire  Queue_10_covMap_write_en; // @[Coverage map for Queue_10]
  reg [29:0] Queue_10_covSum; // @[Sum of coverage map]
  wire  maybe_full_shl;
  wire  maybe_full_pad;
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_cache_io_deq_bits_MPORT_en = 1'h1;
  assign ram_cache_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_cache_io_deq_bits_MPORT_data = ram_cache[ram_cache_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_cache_MPORT_data = io_enq_bits_cache;
  assign ram_cache_MPORT_addr = 1'h0;
  assign ram_cache_MPORT_mask = 1'h1;
  assign ram_cache_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_prot_io_deq_bits_MPORT_en = 1'h1;
  assign ram_prot_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_prot_io_deq_bits_MPORT_data = ram_prot[ram_prot_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_prot_MPORT_data = io_enq_bits_prot;
  assign ram_prot_MPORT_addr = 1'h0;
  assign ram_prot_MPORT_mask = 1'h1;
  assign ram_prot_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign ram_echo_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_extra_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_extra_id_io_deq_bits_MPORT_data = ram_echo_extra_id[ram_echo_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_echo_extra_id_MPORT_data = io_enq_bits_echo_extra_id;
  assign ram_echo_extra_id_MPORT_addr = 1'h0;
  assign ram_echo_extra_id_MPORT_mask = 1'h1;
  assign ram_echo_extra_id_MPORT_en = empty ? _GEN_18 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_burst = empty ? io_enq_bits_burst : ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_cache = empty ? io_enq_bits_cache : ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_prot = empty ? io_enq_bits_prot : ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_echo_extra_id = empty ? io_enq_bits_echo_extra_id : ram_echo_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign Queue_10_covMap_read_en = 1'h1;
  assign Queue_10_covMap_read_addr = Queue_10_covState;
  assign Queue_10_covMap_read_data = Queue_10_covMap[Queue_10_covMap_read_addr]; // @[Coverage map for Queue_10]
  assign Queue_10_covMap_write_data = 1'h1;
  assign Queue_10_covMap_write_addr = Queue_10_covState;
  assign Queue_10_covMap_write_mask = 1'h1;
  assign Queue_10_covMap_write_en = ~metaReset;
  assign maybe_full_shl = maybe_full;
  assign maybe_full_pad = maybe_full_shl;
  assign io_covSum = Queue_10_covSum;
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_cache_MPORT_en & ram_cache_MPORT_mask) begin
      ram_cache[ram_cache_MPORT_addr] <= ram_cache_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_prot_MPORT_en & ram_prot_MPORT_mask) begin
      ram_prot[ram_prot_MPORT_addr] <= ram_prot_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_echo_extra_id_MPORT_en & ram_echo_extra_id_MPORT_mask) begin
      ram_echo_extra_id[ram_echo_extra_id_MPORT_addr] <= ram_echo_extra_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
    Queue_10_covState <= maybe_full_pad;
    if (Queue_10_covMap_write_en & Queue_10_covMap_write_mask) begin
      Queue_10_covMap[Queue_10_covMap_write_addr] <= Queue_10_covMap_write_data; // @[Coverage map for Queue_10]
    end
    if (!(Queue_10_covMap_read_data | metaReset)) begin
      Queue_10_covSum <= Queue_10_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_echo_extra_id[initvar] = _RAND_7[6:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Queue_10_covMap[initvar] = 0; //_10[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  Queue_10_covState = 0; //_9[0:0];
  _RAND_11 = {1{`RANDOM}};
  Queue_10_covSum = 0; //_11[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_12(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input  [7:0]  io_enq_bits_strb,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_strb,
  output        io_deq_bits_last,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_strb [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_strb_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_strb_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_strb_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_strb_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_strb_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_last [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_11 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_11 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  reg  Queue_12_covState; // @[Register tracking Queue_12 state]
  reg  Queue_12_covMap [0:1]; // @[Coverage map for Queue_12]
  wire  Queue_12_covMap_read_en; // @[Coverage map for Queue_12]
  wire  Queue_12_covMap_read_addr; // @[Coverage map for Queue_12]
  wire  Queue_12_covMap_read_data; // @[Coverage map for Queue_12]
  wire  Queue_12_covMap_write_data; // @[Coverage map for Queue_12]
  wire  Queue_12_covMap_write_addr; // @[Coverage map for Queue_12]
  wire  Queue_12_covMap_write_mask; // @[Coverage map for Queue_12]
  wire  Queue_12_covMap_write_en; // @[Coverage map for Queue_12]
  reg [29:0] Queue_12_covSum; // @[Sum of coverage map]
  wire  maybe_full_shl;
  wire  maybe_full_pad;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = 1'h0;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_11 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_strb = empty ? io_enq_bits_strb : ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_last = empty ? io_enq_bits_last : ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign Queue_12_covMap_read_en = 1'h1;
  assign Queue_12_covMap_read_addr = Queue_12_covState;
  assign Queue_12_covMap_read_data = Queue_12_covMap[Queue_12_covMap_read_addr]; // @[Coverage map for Queue_12]
  assign Queue_12_covMap_write_data = 1'h1;
  assign Queue_12_covMap_write_addr = Queue_12_covState;
  assign Queue_12_covMap_write_mask = 1'h1;
  assign Queue_12_covMap_write_en = ~metaReset;
  assign maybe_full_shl = maybe_full;
  assign maybe_full_pad = maybe_full_shl;
  assign io_covSum = Queue_12_covSum;
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
    Queue_12_covState <= maybe_full_pad;
    if (Queue_12_covMap_write_en & Queue_12_covMap_write_mask) begin
      Queue_12_covMap[Queue_12_covMap_write_addr] <= Queue_12_covMap_write_data; // @[Coverage map for Queue_12]
    end
    if (!(Queue_12_covMap_read_data | metaReset)) begin
      Queue_12_covSum <= Queue_12_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_2[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Queue_12_covMap[initvar] = 0; //_5[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  Queue_12_covState = 0; //_4[0:0];
  _RAND_6 = {1{`RANDOM}};
  Queue_12_covSum = 0; //_6[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4Fragmenter(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [6:0]  auto_in_aw_bits_echo_extra_id,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [6:0]  auto_in_b_bits_echo_extra_id,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [6:0]  auto_in_ar_bits_echo_extra_id,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [6:0]  auto_in_r_bits_echo_extra_id,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [6:0]  auto_out_aw_bits_echo_extra_id,
  output        auto_out_aw_bits_echo_real_last,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [6:0]  auto_out_b_bits_echo_extra_id,
  input         auto_out_b_bits_echo_real_last,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [6:0]  auto_out_ar_bits_echo_extra_id,
  output        auto_out_ar_bits_echo_real_last,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [6:0]  auto_out_r_bits_echo_extra_id,
  input         auto_out_r_bits_echo_real_last,
  input         auto_out_r_bits_last,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  deq_clock; // @[Decoupled.scala 361:21]
  wire  deq_reset; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] deq_io_enq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] deq_io_enq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] deq_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] deq_io_enq_bits_burst; // @[Decoupled.scala 361:21]
  wire [3:0] deq_io_enq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] deq_io_enq_bits_prot; // @[Decoupled.scala 361:21]
  wire [6:0] deq_io_enq_bits_echo_extra_id; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] deq_io_deq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] deq_io_deq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] deq_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] deq_io_deq_bits_burst; // @[Decoupled.scala 361:21]
  wire [3:0] deq_io_deq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] deq_io_deq_bits_prot; // @[Decoupled.scala 361:21]
  wire [6:0] deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 361:21]
  wire [29:0] deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  deq_metaReset; // @[Decoupled.scala 361:21]
  wire  deq_1_clock; // @[Decoupled.scala 361:21]
  wire  deq_1_reset; // @[Decoupled.scala 361:21]
  wire  deq_1_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  deq_1_io_enq_valid; // @[Decoupled.scala 361:21]
  wire  deq_1_io_enq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] deq_1_io_enq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] deq_1_io_enq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] deq_1_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] deq_1_io_enq_bits_burst; // @[Decoupled.scala 361:21]
  wire [3:0] deq_1_io_enq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] deq_1_io_enq_bits_prot; // @[Decoupled.scala 361:21]
  wire [6:0] deq_1_io_enq_bits_echo_extra_id; // @[Decoupled.scala 361:21]
  wire  deq_1_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  deq_1_io_deq_valid; // @[Decoupled.scala 361:21]
  wire  deq_1_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] deq_1_io_deq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] deq_1_io_deq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] deq_1_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] deq_1_io_deq_bits_burst; // @[Decoupled.scala 361:21]
  wire [3:0] deq_1_io_deq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] deq_1_io_deq_bits_prot; // @[Decoupled.scala 361:21]
  wire [6:0] deq_1_io_deq_bits_echo_extra_id; // @[Decoupled.scala 361:21]
  wire [29:0] deq_1_io_covSum; // @[Decoupled.scala 361:21]
  wire  deq_1_metaReset; // @[Decoupled.scala 361:21]
  wire  in_w_deq_clock; // @[Decoupled.scala 361:21]
  wire  in_w_deq_reset; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [63:0] in_w_deq_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] in_w_deq_io_enq_bits_strb; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_enq_bits_last; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [63:0] in_w_deq_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] in_w_deq_io_deq_bits_strb; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_deq_bits_last; // @[Decoupled.scala 361:21]
  wire [29:0] in_w_deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  in_w_deq_metaReset; // @[Decoupled.scala 361:21]
  reg  busy; // @[Fragmenter.scala 60:29]
  reg [31:0] r_addr; // @[Fragmenter.scala 61:25]
  reg [7:0] r_len; // @[Fragmenter.scala 62:25]
  wire [7:0] irr_bits_len = deq_io_deq_bits_len; // @[Decoupled.scala 401:19 402:14]
  wire [7:0] len = busy ? r_len : irr_bits_len; // @[Fragmenter.scala 64:23]
  wire [31:0] irr_bits_addr = deq_io_deq_bits_addr; // @[Decoupled.scala 401:19 402:14]
  wire [31:0] addr = busy ? r_addr : irr_bits_addr; // @[Fragmenter.scala 65:23]
  wire [7:0] alignment = addr[10:3]; // @[Fragmenter.scala 69:29]
  wire [31:0] _support1_T = addr ^ 32'h2000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_1 = {1'b0,$signed(_support1_T)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_3 = $signed(_support1_T_1) & 33'sh86032000; // @[Parameters.scala 137:52]
  wire  _support1_T_4 = $signed(_support1_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire [32:0] _support1_T_6 = {1'b0,$signed(addr)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_8 = $signed(_support1_T_6) & 33'sh86012000; // @[Parameters.scala 137:52]
  wire  _support1_T_9 = $signed(_support1_T_8) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_10 = addr ^ 32'h10000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_11 = {1'b0,$signed(_support1_T_10)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_13 = $signed(_support1_T_11) & 33'sh86030000; // @[Parameters.scala 137:52]
  wire  _support1_T_14 = $signed(_support1_T_13) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_15 = addr ^ 32'h2000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_16 = {1'b0,$signed(_support1_T_15)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_18 = $signed(_support1_T_16) & 33'sh86030000; // @[Parameters.scala 137:52]
  wire  _support1_T_19 = $signed(_support1_T_18) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_20 = addr ^ 32'h4000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_21 = {1'b0,$signed(_support1_T_20)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_23 = $signed(_support1_T_21) & 33'sh84000000; // @[Parameters.scala 137:52]
  wire  _support1_T_24 = $signed(_support1_T_23) == 33'sh0; // @[Parameters.scala 137:67]
  wire [32:0] _support1_T_28 = $signed(_support1_T_21) & 33'sh86032000; // @[Parameters.scala 137:52]
  wire  _support1_T_29 = $signed(_support1_T_28) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_30 = addr ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_31 = {1'b0,$signed(_support1_T_30)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_33 = $signed(_support1_T_31) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  _support1_T_34 = $signed(_support1_T_33) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _support1_T_39 = _support1_T_9 | _support1_T_14 | _support1_T_19 | _support1_T_24 | _support1_T_29 |
    _support1_T_34; // @[Fragmenter.scala 76:100]
  wire [7:0] _support1_T_40 = _support1_T_4 ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [2:0] _support1_T_41 = _support1_T_39 ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [7:0] _GEN_16 = {{5'd0}, _support1_T_41}; // @[Mux.scala 27:73]
  wire [7:0] support1 = _support1_T_40 | _GEN_16; // @[Mux.scala 27:73]
  wire [7:0] _GEN_17 = {{1'd0}, len[7:1]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_1 = len | _GEN_17; // @[package.scala 253:43]
  wire [7:0] _GEN_18 = {{2'd0}, _fillLow_T_1[7:2]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_3 = _fillLow_T_1 | _GEN_18; // @[package.scala 253:43]
  wire [7:0] _GEN_19 = {{4'd0}, _fillLow_T_3[7:4]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_5 = _fillLow_T_3 | _GEN_19; // @[package.scala 253:43]
  wire [6:0] fillLow = _fillLow_T_5[7:1]; // @[Fragmenter.scala 85:37]
  wire [7:0] _wipeHigh_T = ~len; // @[Fragmenter.scala 86:32]
  wire [8:0] _wipeHigh_T_1 = {_wipeHigh_T, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_3 = _wipeHigh_T | _wipeHigh_T_1[7:0]; // @[package.scala 244:43]
  wire [9:0] _wipeHigh_T_4 = {_wipeHigh_T_3, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_6 = _wipeHigh_T_3 | _wipeHigh_T_4[7:0]; // @[package.scala 244:43]
  wire [11:0] _wipeHigh_T_7 = {_wipeHigh_T_6, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_9 = _wipeHigh_T_6 | _wipeHigh_T_7[7:0]; // @[package.scala 244:43]
  wire [7:0] wipeHigh = ~_wipeHigh_T_9; // @[Fragmenter.scala 86:24]
  wire [7:0] _GEN_20 = {{1'd0}, fillLow}; // @[Fragmenter.scala 87:32]
  wire [7:0] remain1 = _GEN_20 | wipeHigh; // @[Fragmenter.scala 87:32]
  wire [8:0] _align1_T = {alignment, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_2 = alignment | _align1_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _align1_T_3 = {_align1_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_5 = _align1_T_2 | _align1_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _align1_T_6 = {_align1_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_8 = _align1_T_5 | _align1_T_6[7:0]; // @[package.scala 244:43]
  wire [7:0] align1 = ~_align1_T_8; // @[Fragmenter.scala 88:24]
  wire [7:0] _maxSupported1_T = remain1 & align1; // @[Fragmenter.scala 89:37]
  wire [7:0] maxSupported1 = _maxSupported1_T & support1; // @[Fragmenter.scala 89:46]
  wire [1:0] irr_bits_burst = deq_io_deq_bits_burst; // @[Decoupled.scala 401:19 402:14]
  wire  fixed = irr_bits_burst == 2'h0; // @[Fragmenter.scala 92:34]
  wire [2:0] irr_bits_size = deq_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  wire  narrow = irr_bits_size != 3'h3; // @[Fragmenter.scala 93:34]
  wire  bad = fixed | narrow; // @[Fragmenter.scala 94:25]
  wire [7:0] beats1 = bad ? 8'h0 : maxSupported1; // @[Fragmenter.scala 97:25]
  wire [8:0] _beats_T = {beats1, 1'h0}; // @[package.scala 232:35]
  wire [8:0] _beats_T_1 = _beats_T | 9'h1; // @[package.scala 232:40]
  wire [8:0] _beats_T_2 = {1'h0,beats1}; // @[Cat.scala 31:58]
  wire [8:0] _beats_T_3 = ~_beats_T_2; // @[package.scala 232:53]
  wire [8:0] beats = _beats_T_1 & _beats_T_3; // @[package.scala 232:51]
  wire [15:0] _GEN_39 = {{7'd0}, beats}; // @[Fragmenter.scala 100:38]
  wire [15:0] _inc_addr_T = _GEN_39 << irr_bits_size; // @[Fragmenter.scala 100:38]
  wire [31:0] _GEN_21 = {{16'd0}, _inc_addr_T}; // @[Fragmenter.scala 100:29]
  wire [31:0] inc_addr = addr + _GEN_21; // @[Fragmenter.scala 100:29]
  wire [15:0] _wrapMask_T = {irr_bits_len,8'hff}; // @[Cat.scala 31:58]
  wire [22:0] _GEN_40 = {{7'd0}, _wrapMask_T}; // @[Bundles.scala 31:21]
  wire [22:0] _wrapMask_T_1 = _GEN_40 << irr_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] wrapMask = _wrapMask_T_1[22:8]; // @[Bundles.scala 31:30]
  wire [31:0] _GEN_22 = {{17'd0}, wrapMask}; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T = inc_addr & _GEN_22; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T_1 = ~irr_bits_addr; // @[Fragmenter.scala 104:49]
  wire [31:0] _mux_addr_T_2 = _mux_addr_T_1 | _GEN_22; // @[Fragmenter.scala 104:62]
  wire [31:0] _mux_addr_T_3 = ~_mux_addr_T_2; // @[Fragmenter.scala 104:47]
  wire [31:0] _mux_addr_T_4 = _mux_addr_T | _mux_addr_T_3; // @[Fragmenter.scala 104:45]
  wire  ar_last = beats1 == len; // @[Fragmenter.scala 110:27]
  wire [31:0] _out_bits_addr_T = ~addr; // @[Fragmenter.scala 122:28]
  wire [9:0] _out_bits_addr_T_2 = 10'h7 << irr_bits_size; // @[package.scala 234:77]
  wire [2:0] _out_bits_addr_T_4 = ~_out_bits_addr_T_2[2:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_24 = {{29'd0}, _out_bits_addr_T_4}; // @[Fragmenter.scala 122:34]
  wire [31:0] _out_bits_addr_T_5 = _out_bits_addr_T | _GEN_24; // @[Fragmenter.scala 122:34]
  wire  irr_valid = deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  wire  _T_2 = auto_out_ar_ready & irr_valid; // @[Decoupled.scala 50:35]
  wire [8:0] _GEN_25 = {{1'd0}, len}; // @[Fragmenter.scala 127:25]
  wire [8:0] _r_len_T_1 = _GEN_25 - beats; // @[Fragmenter.scala 127:25]
  wire [8:0] _GEN_4 = _T_2 ? _r_len_T_1 : {{1'd0}, r_len}; // @[Fragmenter.scala 124:27 127:18 62:25]
  reg  busy_1; // @[Fragmenter.scala 60:29]
  reg [31:0] r_addr_1; // @[Fragmenter.scala 61:25]
  reg [7:0] r_len_1; // @[Fragmenter.scala 62:25]
  wire [7:0] irr_1_bits_len = deq_1_io_deq_bits_len; // @[Decoupled.scala 401:19 402:14]
  wire [7:0] len_1 = busy_1 ? r_len_1 : irr_1_bits_len; // @[Fragmenter.scala 64:23]
  wire [31:0] irr_1_bits_addr = deq_1_io_deq_bits_addr; // @[Decoupled.scala 401:19 402:14]
  wire [31:0] addr_1 = busy_1 ? r_addr_1 : irr_1_bits_addr; // @[Fragmenter.scala 65:23]
  wire [7:0] alignment_1 = addr_1[10:3]; // @[Fragmenter.scala 69:29]
  wire [31:0] _support1_T_43 = addr_1 ^ 32'h2000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_44 = {1'b0,$signed(_support1_T_43)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_46 = $signed(_support1_T_44) & 33'sh86002000; // @[Parameters.scala 137:52]
  wire  _support1_T_47 = $signed(_support1_T_46) == 33'sh0; // @[Parameters.scala 137:67]
  wire [32:0] _support1_T_49 = {1'b0,$signed(addr_1)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_51 = $signed(_support1_T_49) & 33'sh82002000; // @[Parameters.scala 137:52]
  wire  _support1_T_52 = $signed(_support1_T_51) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_53 = addr_1 ^ 32'h2000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_54 = {1'b0,$signed(_support1_T_53)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_56 = $signed(_support1_T_54) & 33'sh86000000; // @[Parameters.scala 137:52]
  wire  _support1_T_57 = $signed(_support1_T_56) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_58 = addr_1 ^ 32'h4000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_59 = {1'b0,$signed(_support1_T_58)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_61 = $signed(_support1_T_59) & 33'sh84000000; // @[Parameters.scala 137:52]
  wire  _support1_T_62 = $signed(_support1_T_61) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_63 = addr_1 ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_64 = {1'b0,$signed(_support1_T_63)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_66 = $signed(_support1_T_64) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  _support1_T_67 = $signed(_support1_T_66) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _support1_T_70 = _support1_T_52 | _support1_T_57 | _support1_T_62 | _support1_T_67; // @[Fragmenter.scala 76:100]
  wire [7:0] _support1_T_71 = _support1_T_47 ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [2:0] _support1_T_72 = _support1_T_70 ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [7:0] _GEN_26 = {{5'd0}, _support1_T_72}; // @[Mux.scala 27:73]
  wire [7:0] support1_1 = _support1_T_71 | _GEN_26; // @[Mux.scala 27:73]
  wire [7:0] _GEN_27 = {{1'd0}, len_1[7:1]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_8 = len_1 | _GEN_27; // @[package.scala 253:43]
  wire [7:0] _GEN_28 = {{2'd0}, _fillLow_T_8[7:2]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_10 = _fillLow_T_8 | _GEN_28; // @[package.scala 253:43]
  wire [7:0] _GEN_29 = {{4'd0}, _fillLow_T_10[7:4]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_12 = _fillLow_T_10 | _GEN_29; // @[package.scala 253:43]
  wire [6:0] fillLow_1 = _fillLow_T_12[7:1]; // @[Fragmenter.scala 85:37]
  wire [7:0] _wipeHigh_T_11 = ~len_1; // @[Fragmenter.scala 86:32]
  wire [8:0] _wipeHigh_T_12 = {_wipeHigh_T_11, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_14 = _wipeHigh_T_11 | _wipeHigh_T_12[7:0]; // @[package.scala 244:43]
  wire [9:0] _wipeHigh_T_15 = {_wipeHigh_T_14, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_17 = _wipeHigh_T_14 | _wipeHigh_T_15[7:0]; // @[package.scala 244:43]
  wire [11:0] _wipeHigh_T_18 = {_wipeHigh_T_17, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_20 = _wipeHigh_T_17 | _wipeHigh_T_18[7:0]; // @[package.scala 244:43]
  wire [7:0] wipeHigh_1 = ~_wipeHigh_T_20; // @[Fragmenter.scala 86:24]
  wire [7:0] _GEN_30 = {{1'd0}, fillLow_1}; // @[Fragmenter.scala 87:32]
  wire [7:0] remain1_1 = _GEN_30 | wipeHigh_1; // @[Fragmenter.scala 87:32]
  wire [8:0] _align1_T_10 = {alignment_1, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_12 = alignment_1 | _align1_T_10[7:0]; // @[package.scala 244:43]
  wire [9:0] _align1_T_13 = {_align1_T_12, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_15 = _align1_T_12 | _align1_T_13[7:0]; // @[package.scala 244:43]
  wire [11:0] _align1_T_16 = {_align1_T_15, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_18 = _align1_T_15 | _align1_T_16[7:0]; // @[package.scala 244:43]
  wire [7:0] align1_1 = ~_align1_T_18; // @[Fragmenter.scala 88:24]
  wire [7:0] _maxSupported1_T_1 = remain1_1 & align1_1; // @[Fragmenter.scala 89:37]
  wire [7:0] maxSupported1_1 = _maxSupported1_T_1 & support1_1; // @[Fragmenter.scala 89:46]
  wire [1:0] irr_1_bits_burst = deq_1_io_deq_bits_burst; // @[Decoupled.scala 401:19 402:14]
  wire  fixed_1 = irr_1_bits_burst == 2'h0; // @[Fragmenter.scala 92:34]
  wire [2:0] irr_1_bits_size = deq_1_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  wire  narrow_1 = irr_1_bits_size != 3'h3; // @[Fragmenter.scala 93:34]
  wire  bad_1 = fixed_1 | narrow_1; // @[Fragmenter.scala 94:25]
  wire [7:0] beats1_1 = bad_1 ? 8'h0 : maxSupported1_1; // @[Fragmenter.scala 97:25]
  wire [8:0] _beats_T_4 = {beats1_1, 1'h0}; // @[package.scala 232:35]
  wire [8:0] _beats_T_5 = _beats_T_4 | 9'h1; // @[package.scala 232:40]
  wire [8:0] _beats_T_6 = {1'h0,beats1_1}; // @[Cat.scala 31:58]
  wire [8:0] _beats_T_7 = ~_beats_T_6; // @[package.scala 232:53]
  wire [8:0] w_beats = _beats_T_5 & _beats_T_7; // @[package.scala 232:51]
  wire [15:0] _GEN_56 = {{7'd0}, w_beats}; // @[Fragmenter.scala 100:38]
  wire [15:0] _inc_addr_T_2 = _GEN_56 << irr_1_bits_size; // @[Fragmenter.scala 100:38]
  wire [31:0] _GEN_31 = {{16'd0}, _inc_addr_T_2}; // @[Fragmenter.scala 100:29]
  wire [31:0] inc_addr_1 = addr_1 + _GEN_31; // @[Fragmenter.scala 100:29]
  wire [15:0] _wrapMask_T_2 = {irr_1_bits_len,8'hff}; // @[Cat.scala 31:58]
  wire [22:0] _GEN_57 = {{7'd0}, _wrapMask_T_2}; // @[Bundles.scala 31:21]
  wire [22:0] _wrapMask_T_3 = _GEN_57 << irr_1_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] wrapMask_1 = _wrapMask_T_3[22:8]; // @[Bundles.scala 31:30]
  wire [31:0] _GEN_32 = {{17'd0}, wrapMask_1}; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T_5 = inc_addr_1 & _GEN_32; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T_6 = ~irr_1_bits_addr; // @[Fragmenter.scala 104:49]
  wire [31:0] _mux_addr_T_7 = _mux_addr_T_6 | _GEN_32; // @[Fragmenter.scala 104:62]
  wire [31:0] _mux_addr_T_8 = ~_mux_addr_T_7; // @[Fragmenter.scala 104:47]
  wire [31:0] _mux_addr_T_9 = _mux_addr_T_5 | _mux_addr_T_8; // @[Fragmenter.scala 104:45]
  wire  aw_last = beats1_1 == len_1; // @[Fragmenter.scala 110:27]
  reg [8:0] w_counter; // @[Fragmenter.scala 164:30]
  wire  w_idle = w_counter == 9'h0; // @[Fragmenter.scala 165:30]
  reg  wbeats_latched; // @[Fragmenter.scala 150:35]
  wire  _in_aw_ready_T = w_idle | wbeats_latched; // @[Fragmenter.scala 158:52]
  wire  in_aw_ready = auto_out_aw_ready & (w_idle | wbeats_latched); // @[Fragmenter.scala 158:35]
  wire [31:0] _out_bits_addr_T_7 = ~addr_1; // @[Fragmenter.scala 122:28]
  wire [9:0] _out_bits_addr_T_9 = 10'h7 << irr_1_bits_size; // @[package.scala 234:77]
  wire [2:0] _out_bits_addr_T_11 = ~_out_bits_addr_T_9[2:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_34 = {{29'd0}, _out_bits_addr_T_11}; // @[Fragmenter.scala 122:34]
  wire [31:0] _out_bits_addr_T_12 = _out_bits_addr_T_7 | _GEN_34; // @[Fragmenter.scala 122:34]
  wire  irr_1_valid = deq_1_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  wire  _T_5 = in_aw_ready & irr_1_valid; // @[Decoupled.scala 50:35]
  wire [8:0] _GEN_35 = {{1'd0}, len_1}; // @[Fragmenter.scala 127:25]
  wire [8:0] _r_len_T_3 = _GEN_35 - w_beats; // @[Fragmenter.scala 127:25]
  wire [8:0] _GEN_9 = _T_5 ? _r_len_T_3 : {{1'd0}, r_len_1}; // @[Fragmenter.scala 124:27 127:18 62:25]
  wire  wbeats_valid = irr_1_valid & ~wbeats_latched; // @[Fragmenter.scala 159:35]
  wire  _GEN_10 = wbeats_valid & w_idle | wbeats_latched; // @[Fragmenter.scala 150:35 153:{43,60}]
  wire  bundleOut_0_aw_valid = irr_1_valid & _in_aw_ready_T; // @[Fragmenter.scala 157:35]
  wire  _T_7 = auto_out_aw_ready & bundleOut_0_aw_valid; // @[Decoupled.scala 50:35]
  wire [8:0] _w_todo_T = wbeats_valid ? w_beats : 9'h0; // @[Fragmenter.scala 166:35]
  wire [8:0] w_todo = w_idle ? _w_todo_T : w_counter; // @[Fragmenter.scala 166:23]
  wire  w_last = w_todo == 9'h1; // @[Fragmenter.scala 167:27]
  wire  in_w_valid = in_w_deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  wire  _bundleOut_0_w_valid_T_1 = ~w_idle | wbeats_valid; // @[Fragmenter.scala 173:51]
  wire  bundleOut_0_w_valid = in_w_valid & (~w_idle | wbeats_valid); // @[Fragmenter.scala 173:33]
  wire  _w_counter_T = auto_out_w_ready & bundleOut_0_w_valid; // @[Decoupled.scala 50:35]
  wire [8:0] _GEN_36 = {{8'd0}, _w_counter_T}; // @[Fragmenter.scala 168:27]
  wire [8:0] _w_counter_T_2 = w_todo - _GEN_36; // @[Fragmenter.scala 168:27]
  wire  _T_13 = ~reset; // @[Fragmenter.scala 169:14]
  wire  in_w_bits_last = in_w_deq_io_deq_bits_last; // @[Decoupled.scala 401:19 402:14]
  wire  bundleOut_0_b_ready = auto_in_b_ready | ~auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 189:33]
  reg [1:0] error_0; // @[Fragmenter.scala 192:26]
  reg [1:0] error_1; // @[Fragmenter.scala 192:26]
  wire [1:0] _GEN_13 = auto_out_b_bits_id ? error_1 : error_0; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _T_22 = 2'h1 << auto_out_b_bits_id; // @[OneHot.scala 64:12]
  wire  _T_26 = bundleOut_0_b_ready & auto_out_b_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _error_0_T = error_0 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_1_T = error_1 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  reg [6:0] AXI4Fragmenter_covState; // @[Register tracking AXI4Fragmenter state]
  reg  AXI4Fragmenter_covMap [0:127]; // @[Coverage map for AXI4Fragmenter]
  wire  AXI4Fragmenter_covMap_read_en; // @[Coverage map for AXI4Fragmenter]
  wire [6:0] AXI4Fragmenter_covMap_read_addr; // @[Coverage map for AXI4Fragmenter]
  wire  AXI4Fragmenter_covMap_read_data; // @[Coverage map for AXI4Fragmenter]
  wire  AXI4Fragmenter_covMap_write_data; // @[Coverage map for AXI4Fragmenter]
  wire [6:0] AXI4Fragmenter_covMap_write_addr; // @[Coverage map for AXI4Fragmenter]
  wire  AXI4Fragmenter_covMap_write_mask; // @[Coverage map for AXI4Fragmenter]
  wire  AXI4Fragmenter_covMap_write_en; // @[Coverage map for AXI4Fragmenter]
  reg [29:0] AXI4Fragmenter_covSum; // @[Sum of coverage map]
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  busy_shl;
  wire [6:0] busy_pad;
  wire [1:0] wbeats_latched_shl;
  wire [6:0] wbeats_latched_pad;
  wire [2:0] busy_1_shl;
  wire [6:0] busy_1_pad;
  wire [3:0] mux_cond_0_shl;
  wire [6:0] mux_cond_0_pad;
  wire [4:0] mux_cond_1_shl;
  wire [6:0] mux_cond_1_pad;
  wire [5:0] mux_cond_2_shl;
  wire [6:0] mux_cond_2_pad;
  wire [6:0] mux_cond_3_shl;
  wire [6:0] mux_cond_3_pad;
  wire [6:0] AXI4Fragmenter_xor4;
  wire [6:0] AXI4Fragmenter_xor1;
  wire [6:0] AXI4Fragmenter_xor5;
  wire [6:0] AXI4Fragmenter_xor6;
  wire [6:0] AXI4Fragmenter_xor2;
  wire [6:0] AXI4Fragmenter_xor0;
  wire [29:0] deq_sum;
  wire [29:0] deq_1_sum;
  wire [29:0] in_w_deq_sum;
  Queue_10 deq ( // @[Decoupled.scala 361:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_id(deq_io_enq_bits_id),
    .io_enq_bits_addr(deq_io_enq_bits_addr),
    .io_enq_bits_len(deq_io_enq_bits_len),
    .io_enq_bits_size(deq_io_enq_bits_size),
    .io_enq_bits_burst(deq_io_enq_bits_burst),
    .io_enq_bits_cache(deq_io_enq_bits_cache),
    .io_enq_bits_prot(deq_io_enq_bits_prot),
    .io_enq_bits_echo_extra_id(deq_io_enq_bits_echo_extra_id),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_id(deq_io_deq_bits_id),
    .io_deq_bits_addr(deq_io_deq_bits_addr),
    .io_deq_bits_len(deq_io_deq_bits_len),
    .io_deq_bits_size(deq_io_deq_bits_size),
    .io_deq_bits_burst(deq_io_deq_bits_burst),
    .io_deq_bits_cache(deq_io_deq_bits_cache),
    .io_deq_bits_prot(deq_io_deq_bits_prot),
    .io_deq_bits_echo_extra_id(deq_io_deq_bits_echo_extra_id),
    .io_covSum(deq_io_covSum),
    .metaReset(deq_metaReset)
  );
  Queue_10 deq_1 ( // @[Decoupled.scala 361:21]
    .clock(deq_1_clock),
    .reset(deq_1_reset),
    .io_enq_ready(deq_1_io_enq_ready),
    .io_enq_valid(deq_1_io_enq_valid),
    .io_enq_bits_id(deq_1_io_enq_bits_id),
    .io_enq_bits_addr(deq_1_io_enq_bits_addr),
    .io_enq_bits_len(deq_1_io_enq_bits_len),
    .io_enq_bits_size(deq_1_io_enq_bits_size),
    .io_enq_bits_burst(deq_1_io_enq_bits_burst),
    .io_enq_bits_cache(deq_1_io_enq_bits_cache),
    .io_enq_bits_prot(deq_1_io_enq_bits_prot),
    .io_enq_bits_echo_extra_id(deq_1_io_enq_bits_echo_extra_id),
    .io_deq_ready(deq_1_io_deq_ready),
    .io_deq_valid(deq_1_io_deq_valid),
    .io_deq_bits_id(deq_1_io_deq_bits_id),
    .io_deq_bits_addr(deq_1_io_deq_bits_addr),
    .io_deq_bits_len(deq_1_io_deq_bits_len),
    .io_deq_bits_size(deq_1_io_deq_bits_size),
    .io_deq_bits_burst(deq_1_io_deq_bits_burst),
    .io_deq_bits_cache(deq_1_io_deq_bits_cache),
    .io_deq_bits_prot(deq_1_io_deq_bits_prot),
    .io_deq_bits_echo_extra_id(deq_1_io_deq_bits_echo_extra_id),
    .io_covSum(deq_1_io_covSum),
    .metaReset(deq_1_metaReset)
  );
  Queue_12 in_w_deq ( // @[Decoupled.scala 361:21]
    .clock(in_w_deq_clock),
    .reset(in_w_deq_reset),
    .io_enq_ready(in_w_deq_io_enq_ready),
    .io_enq_valid(in_w_deq_io_enq_valid),
    .io_enq_bits_data(in_w_deq_io_enq_bits_data),
    .io_enq_bits_strb(in_w_deq_io_enq_bits_strb),
    .io_enq_bits_last(in_w_deq_io_enq_bits_last),
    .io_deq_ready(in_w_deq_io_deq_ready),
    .io_deq_valid(in_w_deq_io_deq_valid),
    .io_deq_bits_data(in_w_deq_io_deq_bits_data),
    .io_deq_bits_strb(in_w_deq_io_deq_bits_strb),
    .io_deq_bits_last(in_w_deq_io_deq_bits_last),
    .io_covSum(in_w_deq_io_covSum),
    .metaReset(in_w_deq_metaReset)
  );
  assign auto_in_aw_ready = deq_1_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_w_ready = in_w_deq_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_b_valid = auto_out_b_valid & auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 188:33]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp | _GEN_13; // @[Fragmenter.scala 193:41]
  assign auto_in_b_bits_echo_extra_id = auto_out_b_bits_echo_extra_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_ar_ready = deq_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_echo_extra_id = auto_out_r_bits_echo_extra_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last & auto_out_r_bits_echo_real_last; // @[Fragmenter.scala 183:41]
  assign auto_out_aw_valid = irr_1_valid & _in_aw_ready_T; // @[Fragmenter.scala 157:35]
  assign auto_out_aw_bits_id = deq_1_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_addr = ~_out_bits_addr_T_12; // @[Fragmenter.scala 122:26]
  assign auto_out_aw_bits_len = bad_1 ? 8'h0 : maxSupported1_1; // @[Fragmenter.scala 97:25]
  assign auto_out_aw_bits_size = deq_1_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_cache = deq_1_io_deq_bits_cache; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_prot = deq_1_io_deq_bits_prot; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_echo_extra_id = deq_1_io_deq_bits_echo_extra_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_echo_real_last = beats1_1 == len_1; // @[Fragmenter.scala 110:27]
  assign auto_out_w_valid = in_w_valid & (~w_idle | wbeats_valid); // @[Fragmenter.scala 173:33]
  assign auto_out_w_bits_data = in_w_deq_io_deq_bits_data; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_w_bits_strb = in_w_deq_io_deq_bits_strb; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_w_bits_last = w_todo == 9'h1; // @[Fragmenter.scala 167:27]
  assign auto_out_b_ready = auto_in_b_ready | ~auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 189:33]
  assign auto_out_ar_valid = deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  assign auto_out_ar_bits_id = deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_addr = ~_out_bits_addr_T_5; // @[Fragmenter.scala 122:26]
  assign auto_out_ar_bits_len = bad ? 8'h0 : maxSupported1; // @[Fragmenter.scala 97:25]
  assign auto_out_ar_bits_size = deq_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_cache = deq_io_deq_bits_cache; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_prot = deq_io_deq_bits_prot; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_echo_extra_id = deq_io_deq_bits_echo_extra_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_echo_real_last = beats1 == len; // @[Fragmenter.scala 110:27]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = auto_in_ar_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_echo_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_deq_ready = auto_out_ar_ready & ar_last; // @[Fragmenter.scala 111:30]
  assign deq_1_clock = clock;
  assign deq_1_reset = reset;
  assign deq_1_io_enq_valid = auto_in_aw_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_echo_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_deq_ready = in_aw_ready & aw_last; // @[Fragmenter.scala 111:30]
  assign in_w_deq_clock = clock;
  assign in_w_deq_reset = reset;
  assign in_w_deq_io_enq_valid = auto_in_w_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_w_deq_io_enq_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_w_deq_io_enq_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_w_deq_io_enq_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_w_deq_io_deq_ready = auto_out_w_ready & _bundleOut_0_w_valid_T_1; // @[Fragmenter.scala 174:33]
  assign AXI4Fragmenter_covMap_read_en = 1'h1;
  assign AXI4Fragmenter_covMap_read_addr = AXI4Fragmenter_covState;
  assign AXI4Fragmenter_covMap_read_data = AXI4Fragmenter_covMap[AXI4Fragmenter_covMap_read_addr]; // @[Coverage map for AXI4Fragmenter]
  assign AXI4Fragmenter_covMap_write_data = 1'h1;
  assign AXI4Fragmenter_covMap_write_addr = AXI4Fragmenter_covState;
  assign AXI4Fragmenter_covMap_write_mask = 1'h1;
  assign AXI4Fragmenter_covMap_write_en = ~metaReset;
  assign mux_cond_0 = _support1_T_47;
  assign mux_cond_1 = _support1_T_4;
  assign mux_cond_2 = _support1_T_39;
  assign mux_cond_3 = _support1_T_70;
  assign busy_shl = busy;
  assign busy_pad = {6'h0,busy_shl};
  assign wbeats_latched_shl = {wbeats_latched, 1'h0};
  assign wbeats_latched_pad = {5'h0,wbeats_latched_shl};
  assign busy_1_shl = {busy_1, 2'h0};
  assign busy_1_pad = {4'h0,busy_1_shl};
  assign mux_cond_0_shl = {mux_cond_0, 3'h0};
  assign mux_cond_0_pad = {3'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 4'h0};
  assign mux_cond_1_pad = {2'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 5'h0};
  assign mux_cond_2_pad = {1'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 6'h0};
  assign mux_cond_3_pad = mux_cond_3_shl;
  assign AXI4Fragmenter_xor4 = wbeats_latched_pad ^ busy_1_pad;
  assign AXI4Fragmenter_xor1 = busy_pad ^ AXI4Fragmenter_xor4;
  assign AXI4Fragmenter_xor5 = mux_cond_0_pad ^ mux_cond_1_pad;
  assign AXI4Fragmenter_xor6 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign AXI4Fragmenter_xor2 = AXI4Fragmenter_xor5 ^ AXI4Fragmenter_xor6;
  assign AXI4Fragmenter_xor0 = AXI4Fragmenter_xor1 ^ AXI4Fragmenter_xor2;
  assign deq_sum = AXI4Fragmenter_covSum + deq_io_covSum;
  assign deq_1_sum = deq_sum + deq_1_io_covSum;
  assign in_w_deq_sum = deq_1_sum + in_w_deq_io_covSum;
  assign io_covSum = in_w_deq_sum;
  assign deq_metaReset = metaReset;
  assign deq_1_metaReset = metaReset;
  assign in_w_deq_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 60:29]
      busy <= 1'h0; // @[Fragmenter.scala 60:29]
    end else if (_T_2) begin
      busy <= ~ar_last;
    end
    if (_T_2) begin // @[Fragmenter.scala 124:27]
      if (fixed) begin
        r_addr <= irr_bits_addr;
      end else if (irr_bits_burst == 2'h2) begin
        r_addr <= _mux_addr_T_4;
      end else begin
        r_addr <= inc_addr;
      end
    end
    r_len <= _GEN_4[7:0];
    if (reset) begin // @[Fragmenter.scala 60:29]
      busy_1 <= 1'h0; // @[Fragmenter.scala 60:29]
    end else if (_T_5) begin
      busy_1 <= ~aw_last;
    end
    if (_T_5) begin // @[Fragmenter.scala 124:27]
      if (fixed_1) begin
        r_addr_1 <= irr_1_bits_addr;
      end else if (irr_1_bits_burst == 2'h2) begin
        r_addr_1 <= _mux_addr_T_9;
      end else begin
        r_addr_1 <= inc_addr_1;
      end
    end
    r_len_1 <= _GEN_9[7:0];
    if (reset) begin // @[Fragmenter.scala 164:30]
      w_counter <= 9'h0; // @[Fragmenter.scala 164:30]
    end else begin
      w_counter <= _w_counter_T_2; // @[Fragmenter.scala 168:17]
    end
    if (reset) begin // @[Fragmenter.scala 150:35]
      wbeats_latched <= 1'h0; // @[Fragmenter.scala 150:35]
    end else if (_T_7) begin
      wbeats_latched <= 1'h0;
    end else begin
      wbeats_latched <= _GEN_10;
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_0 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[0] & _T_26) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_0 <= 2'h0;
      end else begin
        error_0 <= _error_0_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_1 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[1] & _T_26) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_1 <= 2'h0;
      end else begin
        error_1 <= _error_1_T;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_w_counter_T | w_todo != 9'h0) & ~reset) begin
          $fatal; // @[Fragmenter.scala 169:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~_w_counter_T | w_todo != 9'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:169 assert (!out.w.fire() || w_todo =/= UInt(0)) // underflow impossible\n"
            ); // @[Fragmenter.scala 169:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~bundleOut_0_w_valid | ~in_w_bits_last | w_last) & _T_13) begin
          $fatal; // @[Fragmenter.scala 178:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(~bundleOut_0_w_valid | ~in_w_bits_last | w_last)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:178 assert (!out.w.valid || !in_w.bits.last || w_last)\n"); // @[Fragmenter.scala 178:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    AXI4Fragmenter_covState <= AXI4Fragmenter_xor0;
    if (AXI4Fragmenter_covMap_write_en & AXI4Fragmenter_covMap_write_mask) begin
      AXI4Fragmenter_covMap[AXI4Fragmenter_covMap_write_addr] <= AXI4Fragmenter_covMap_write_data; // @[Coverage map for AXI4Fragmenter]
    end
    if (!(AXI4Fragmenter_covMap_read_data | metaReset)) begin
      AXI4Fragmenter_covSum <= AXI4Fragmenter_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    AXI4Fragmenter_covMap[initvar] = 0; //_11[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_len = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  busy_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_addr_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  r_len_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  w_counter = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  wbeats_latched = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  error_0 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  error_1 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  AXI4Fragmenter_covState = 0; //_10[6:0];
  _RAND_12 = {1{`RANDOM}};
  AXI4Fragmenter_covSum = 0; //_12[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4IdIndexer(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [7:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [7:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [7:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [7:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [6:0]  auto_out_aw_bits_echo_extra_id,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [6:0]  auto_out_b_bits_echo_extra_id,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [6:0]  auto_out_ar_bits_echo_extra_id,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [6:0]  auto_out_r_bits_echo_extra_id,
  input         auto_out_r_bits_last,
  output [29:0] io_covSum
);
  wire [29:0] AXI4IdIndexer_covSum;
  assign auto_in_aw_ready = auto_out_aw_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_id = {auto_out_b_bits_echo_extra_id,auto_out_b_bits_id}; // @[Cat.scala 31:58]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_id = {auto_out_r_bits_echo_extra_id,auto_out_r_bits_id}; // @[Cat.scala 31:58]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id[0]; // @[Nodes.scala 1207:84 BundleMap.scala 247:19]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_echo_extra_id = auto_in_aw_bits_id[7:1]; // @[IdIndexer.scala 71:56]
  assign auto_out_w_valid = auto_in_w_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id[0]; // @[Nodes.scala 1207:84 BundleMap.scala 247:19]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_echo_extra_id = auto_in_ar_bits_id[7:1]; // @[IdIndexer.scala 70:56]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign AXI4IdIndexer_covSum = 30'h0;
  assign io_covSum = AXI4IdIndexer_covSum;
endmodule
module TLInterconnectCoupler_5(
  input         clock,
  input         reset,
  output        auto_axi4index_in_aw_ready,
  input         auto_axi4index_in_aw_valid,
  input  [7:0]  auto_axi4index_in_aw_bits_id,
  input  [31:0] auto_axi4index_in_aw_bits_addr,
  input  [7:0]  auto_axi4index_in_aw_bits_len,
  input  [2:0]  auto_axi4index_in_aw_bits_size,
  input  [1:0]  auto_axi4index_in_aw_bits_burst,
  input  [3:0]  auto_axi4index_in_aw_bits_cache,
  input  [2:0]  auto_axi4index_in_aw_bits_prot,
  output        auto_axi4index_in_w_ready,
  input         auto_axi4index_in_w_valid,
  input  [63:0] auto_axi4index_in_w_bits_data,
  input  [7:0]  auto_axi4index_in_w_bits_strb,
  input         auto_axi4index_in_w_bits_last,
  input         auto_axi4index_in_b_ready,
  output        auto_axi4index_in_b_valid,
  output [7:0]  auto_axi4index_in_b_bits_id,
  output [1:0]  auto_axi4index_in_b_bits_resp,
  output        auto_axi4index_in_ar_ready,
  input         auto_axi4index_in_ar_valid,
  input  [7:0]  auto_axi4index_in_ar_bits_id,
  input  [31:0] auto_axi4index_in_ar_bits_addr,
  input  [7:0]  auto_axi4index_in_ar_bits_len,
  input  [2:0]  auto_axi4index_in_ar_bits_size,
  input  [1:0]  auto_axi4index_in_ar_bits_burst,
  input  [3:0]  auto_axi4index_in_ar_bits_cache,
  input  [2:0]  auto_axi4index_in_ar_bits_prot,
  input         auto_axi4index_in_r_ready,
  output        auto_axi4index_in_r_valid,
  output [7:0]  auto_axi4index_in_r_bits_id,
  output [63:0] auto_axi4index_in_r_bits_data,
  output [1:0]  auto_axi4index_in_r_bits_resp,
  output        auto_axi4index_in_r_bits_last,
  input         auto_tl_out_a_ready,
  output        auto_tl_out_a_valid,
  output [2:0]  auto_tl_out_a_bits_opcode,
  output [2:0]  auto_tl_out_a_bits_param,
  output [3:0]  auto_tl_out_a_bits_size,
  output [3:0]  auto_tl_out_a_bits_source,
  output [31:0] auto_tl_out_a_bits_address,
  output        auto_tl_out_a_bits_user_amba_prot_bufferable,
  output        auto_tl_out_a_bits_user_amba_prot_modifiable,
  output        auto_tl_out_a_bits_user_amba_prot_readalloc,
  output        auto_tl_out_a_bits_user_amba_prot_writealloc,
  output        auto_tl_out_a_bits_user_amba_prot_privileged,
  output        auto_tl_out_a_bits_user_amba_prot_secure,
  output        auto_tl_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_tl_out_a_bits_mask,
  output [63:0] auto_tl_out_a_bits_data,
  output        auto_tl_out_d_ready,
  input         auto_tl_out_d_valid,
  input  [2:0]  auto_tl_out_d_bits_opcode,
  input  [3:0]  auto_tl_out_d_bits_size,
  input  [3:0]  auto_tl_out_d_bits_source,
  input         auto_tl_out_d_bits_denied,
  input  [63:0] auto_tl_out_d_bits_data,
  input         auto_tl_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  buffer_clock; // @[Buffer.scala 68:28]
  wire  buffer_reset; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28]
  wire [31:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_bufferable; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_modifiable; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_readalloc; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_writealloc; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_privileged; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_secure; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_fetch; // @[Buffer.scala 68:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28]
  wire [31:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_bufferable; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_modifiable; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_readalloc; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_writealloc; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_privileged; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_secure; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_fetch; // @[Buffer.scala 68:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire [29:0] buffer_io_covSum; // @[Buffer.scala 68:28]
  wire  fixer_clock; // @[FIFOFixer.scala 144:27]
  wire  fixer_reset; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_in_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_in_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_out_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_out_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire [29:0] fixer_io_covSum; // @[FIFOFixer.scala 144:27]
  wire  fixer_metaReset; // @[FIFOFixer.scala 144:27]
  wire  widget_auto_in_a_ready;
  wire  widget_auto_in_a_valid;
  wire [2:0] widget_auto_in_a_bits_opcode;
  wire [3:0] widget_auto_in_a_bits_size;
  wire [3:0] widget_auto_in_a_bits_source;
  wire [31:0] widget_auto_in_a_bits_address;
  wire  widget_auto_in_a_bits_user_amba_prot_bufferable;
  wire  widget_auto_in_a_bits_user_amba_prot_modifiable;
  wire  widget_auto_in_a_bits_user_amba_prot_readalloc;
  wire  widget_auto_in_a_bits_user_amba_prot_writealloc;
  wire  widget_auto_in_a_bits_user_amba_prot_privileged;
  wire  widget_auto_in_a_bits_user_amba_prot_secure;
  wire  widget_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] widget_auto_in_a_bits_mask;
  wire [63:0] widget_auto_in_a_bits_data;
  wire  widget_auto_in_d_ready;
  wire  widget_auto_in_d_valid;
  wire [2:0] widget_auto_in_d_bits_opcode;
  wire [3:0] widget_auto_in_d_bits_size;
  wire [3:0] widget_auto_in_d_bits_source;
  wire  widget_auto_in_d_bits_denied;
  wire [63:0] widget_auto_in_d_bits_data;
  wire  widget_auto_in_d_bits_corrupt;
  wire  widget_auto_out_a_ready;
  wire  widget_auto_out_a_valid;
  wire [2:0] widget_auto_out_a_bits_opcode;
  wire [3:0] widget_auto_out_a_bits_size;
  wire [3:0] widget_auto_out_a_bits_source;
  wire [31:0] widget_auto_out_a_bits_address;
  wire  widget_auto_out_a_bits_user_amba_prot_bufferable;
  wire  widget_auto_out_a_bits_user_amba_prot_modifiable;
  wire  widget_auto_out_a_bits_user_amba_prot_readalloc;
  wire  widget_auto_out_a_bits_user_amba_prot_writealloc;
  wire  widget_auto_out_a_bits_user_amba_prot_privileged;
  wire  widget_auto_out_a_bits_user_amba_prot_secure;
  wire  widget_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] widget_auto_out_a_bits_mask;
  wire [63:0] widget_auto_out_a_bits_data;
  wire  widget_auto_out_d_ready;
  wire  widget_auto_out_d_valid;
  wire [2:0] widget_auto_out_d_bits_opcode;
  wire [3:0] widget_auto_out_d_bits_size;
  wire [3:0] widget_auto_out_d_bits_source;
  wire  widget_auto_out_d_bits_denied;
  wire [63:0] widget_auto_out_d_bits_data;
  wire  widget_auto_out_d_bits_corrupt;
  wire  axi42tl_clock; // @[ToTL.scala 216:29]
  wire  axi42tl_reset; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_aw_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_aw_valid; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_aw_bits_id; // @[ToTL.scala 216:29]
  wire [31:0] axi42tl_auto_in_aw_bits_addr; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_in_aw_bits_len; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_aw_bits_size; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_in_aw_bits_cache; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_aw_bits_prot; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_w_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_w_valid; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_in_w_bits_data; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_in_w_bits_strb; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_w_bits_last; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_b_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_b_valid; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_b_bits_id; // @[ToTL.scala 216:29]
  wire [1:0] axi42tl_auto_in_b_bits_resp; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_ar_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_ar_valid; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_ar_bits_id; // @[ToTL.scala 216:29]
  wire [31:0] axi42tl_auto_in_ar_bits_addr; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_in_ar_bits_len; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_ar_bits_size; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_in_ar_bits_cache; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_ar_bits_prot; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_r_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_r_valid; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_r_bits_id; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_in_r_bits_data; // @[ToTL.scala 216:29]
  wire [1:0] axi42tl_auto_in_r_bits_resp; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_r_bits_last; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_valid; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_out_a_bits_opcode; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_out_a_bits_size; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_out_a_bits_source; // @[ToTL.scala 216:29]
  wire [31:0] axi42tl_auto_out_a_bits_address; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_bufferable; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_modifiable; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_readalloc; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_writealloc; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_privileged; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_secure; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_fetch; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_out_a_bits_mask; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_out_a_bits_data; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_valid; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_out_d_bits_opcode; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_out_d_bits_size; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_out_d_bits_source; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_bits_denied; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_out_d_bits_data; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_bits_corrupt; // @[ToTL.scala 216:29]
  wire [29:0] axi42tl_io_covSum; // @[ToTL.scala 216:29]
  wire  axi42tl_metaReset; // @[ToTL.scala 216:29]
  wire  axi4yank_clock; // @[UserYanker.scala 105:30]
  wire  axi4yank_reset; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_valid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_in_aw_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_aw_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_aw_bits_size; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_aw_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_aw_bits_prot; // @[UserYanker.scala 105:30]
  wire [6:0] axi4yank_auto_in_aw_bits_echo_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_bits_echo_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_w_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_w_valid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_in_w_bits_data; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_w_bits_strb; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_w_bits_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_b_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_b_valid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_b_bits_id; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_b_bits_resp; // @[UserYanker.scala 105:30]
  wire [6:0] axi4yank_auto_in_b_bits_echo_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_b_bits_echo_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_valid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_in_ar_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_ar_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_ar_bits_size; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_ar_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_ar_bits_prot; // @[UserYanker.scala 105:30]
  wire [6:0] axi4yank_auto_in_ar_bits_echo_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_bits_echo_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_valid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_bits_id; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_in_r_bits_data; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_r_bits_resp; // @[UserYanker.scala 105:30]
  wire [6:0] axi4yank_auto_in_r_bits_echo_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_bits_echo_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_bits_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_aw_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_aw_valid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_aw_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_out_aw_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_aw_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_aw_bits_size; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_aw_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_aw_bits_prot; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_w_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_w_valid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_out_w_bits_data; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_w_bits_strb; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_w_bits_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_b_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_b_valid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_b_bits_id; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_b_bits_resp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_ar_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_ar_valid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_ar_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_out_ar_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_ar_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_ar_bits_size; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_ar_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_ar_bits_prot; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_valid; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_bits_id; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_out_r_bits_data; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_r_bits_resp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_bits_last; // @[UserYanker.scala 105:30]
  wire [29:0] axi4yank_io_covSum; // @[UserYanker.scala 105:30]
  wire  axi4frag_clock; // @[Fragmenter.scala 205:30]
  wire  axi4frag_reset; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_aw_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_aw_valid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_aw_bits_id; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_in_aw_bits_addr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_in_aw_bits_len; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_aw_bits_size; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_aw_bits_burst; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_in_aw_bits_cache; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_aw_bits_prot; // @[Fragmenter.scala 205:30]
  wire [6:0] axi4frag_auto_in_aw_bits_echo_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_w_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_w_valid; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_in_w_bits_data; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_in_w_bits_strb; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_w_bits_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_b_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_b_valid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_b_bits_id; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_b_bits_resp; // @[Fragmenter.scala 205:30]
  wire [6:0] axi4frag_auto_in_b_bits_echo_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_ar_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_ar_valid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_ar_bits_id; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_in_ar_bits_addr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_in_ar_bits_len; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_ar_bits_size; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_ar_bits_burst; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_in_ar_bits_cache; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_ar_bits_prot; // @[Fragmenter.scala 205:30]
  wire [6:0] axi4frag_auto_in_ar_bits_echo_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_r_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_r_valid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_r_bits_id; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_in_r_bits_data; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_r_bits_resp; // @[Fragmenter.scala 205:30]
  wire [6:0] axi4frag_auto_in_r_bits_echo_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_r_bits_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_aw_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_aw_valid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_aw_bits_id; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_out_aw_bits_addr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_out_aw_bits_len; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_aw_bits_size; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_out_aw_bits_cache; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_aw_bits_prot; // @[Fragmenter.scala 205:30]
  wire [6:0] axi4frag_auto_out_aw_bits_echo_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_aw_bits_echo_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_w_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_w_valid; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_out_w_bits_data; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_out_w_bits_strb; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_w_bits_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_b_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_b_valid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_b_bits_id; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_out_b_bits_resp; // @[Fragmenter.scala 205:30]
  wire [6:0] axi4frag_auto_out_b_bits_echo_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_ar_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_ar_valid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_ar_bits_id; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_out_ar_bits_addr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_out_ar_bits_len; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_ar_bits_size; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_out_ar_bits_cache; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_ar_bits_prot; // @[Fragmenter.scala 205:30]
  wire [6:0] axi4frag_auto_out_ar_bits_echo_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_ar_bits_echo_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_r_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_r_valid; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_r_bits_id; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_out_r_bits_data; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_out_r_bits_resp; // @[Fragmenter.scala 205:30]
  wire [6:0] axi4frag_auto_out_r_bits_echo_extra_id; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_r_bits_echo_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_r_bits_last; // @[Fragmenter.scala 205:30]
  wire [29:0] axi4frag_io_covSum; // @[Fragmenter.scala 205:30]
  wire  axi4frag_metaReset; // @[Fragmenter.scala 205:30]
  wire  axi4index_auto_in_aw_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_aw_valid; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_aw_bits_id; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_in_aw_bits_addr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_aw_bits_len; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_aw_bits_size; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_aw_bits_burst; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_aw_bits_cache; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_aw_bits_prot; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_w_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_w_valid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_in_w_bits_data; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_w_bits_strb; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_w_bits_last; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_b_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_b_valid; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_b_bits_id; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_b_bits_resp; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_ar_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_ar_valid; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_ar_bits_id; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_in_ar_bits_addr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_ar_bits_len; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_ar_bits_size; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_ar_bits_burst; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_ar_bits_cache; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_ar_bits_prot; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_r_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_r_valid; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_r_bits_id; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_in_r_bits_data; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_r_bits_resp; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_r_bits_last; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_aw_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_aw_valid; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_aw_bits_id; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_out_aw_bits_addr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_out_aw_bits_len; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_aw_bits_size; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_aw_bits_burst; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_aw_bits_cache; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_aw_bits_prot; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_auto_out_aw_bits_echo_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_w_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_w_valid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_out_w_bits_data; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_out_w_bits_strb; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_w_bits_last; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_b_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_b_valid; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_b_bits_id; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_b_bits_resp; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_auto_out_b_bits_echo_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_ar_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_ar_valid; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_ar_bits_id; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_out_ar_bits_addr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_out_ar_bits_len; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_ar_bits_size; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_ar_bits_burst; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_ar_bits_cache; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_ar_bits_prot; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_auto_out_ar_bits_echo_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_r_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_r_valid; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_r_bits_id; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_out_r_bits_data; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_r_bits_resp; // @[IdIndexer.scala 91:31]
  wire [6:0] axi4index_auto_out_r_bits_echo_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_r_bits_last; // @[IdIndexer.scala 91:31]
  wire [29:0] axi4index_io_covSum; // @[IdIndexer.scala 91:31]
  wire [29:0] TLInterconnectCoupler_5_covSum;
  wire [29:0] fixer_sum;
  wire [29:0] axi42tl_sum;
  wire [29:0] axi4yank_sum;
  wire [29:0] axi4frag_sum;
  wire [29:0] buffer_sum;
  wire [29:0] axi4index_sum;
  TLBuffer_2 buffer ( // @[Buffer.scala 68:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(buffer_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(buffer_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(buffer_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(buffer_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(buffer_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(buffer_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(buffer_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(buffer_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(buffer_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(buffer_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(buffer_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(buffer_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(buffer_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(buffer_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt),
    .io_covSum(buffer_io_covSum)
  );
  TLFIFOFixer_2 fixer ( // @[FIFOFixer.scala 144:27]
    .clock(fixer_clock),
    .reset(fixer_reset),
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(fixer_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(fixer_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(fixer_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(fixer_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(fixer_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(fixer_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(fixer_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_auto_in_a_bits_data),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(fixer_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(fixer_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(fixer_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(fixer_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(fixer_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(fixer_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(fixer_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_auto_out_a_bits_data),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt),
    .io_covSum(fixer_io_covSum),
    .metaReset(fixer_metaReset)
  );
  AXI4ToTL axi42tl ( // @[ToTL.scala 216:29]
    .clock(axi42tl_clock),
    .reset(axi42tl_reset),
    .auto_in_aw_ready(axi42tl_auto_in_aw_ready),
    .auto_in_aw_valid(axi42tl_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi42tl_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi42tl_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi42tl_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi42tl_auto_in_aw_bits_size),
    .auto_in_aw_bits_cache(axi42tl_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi42tl_auto_in_aw_bits_prot),
    .auto_in_w_ready(axi42tl_auto_in_w_ready),
    .auto_in_w_valid(axi42tl_auto_in_w_valid),
    .auto_in_w_bits_data(axi42tl_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi42tl_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi42tl_auto_in_w_bits_last),
    .auto_in_b_ready(axi42tl_auto_in_b_ready),
    .auto_in_b_valid(axi42tl_auto_in_b_valid),
    .auto_in_b_bits_id(axi42tl_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi42tl_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi42tl_auto_in_ar_ready),
    .auto_in_ar_valid(axi42tl_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi42tl_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi42tl_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi42tl_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi42tl_auto_in_ar_bits_size),
    .auto_in_ar_bits_cache(axi42tl_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi42tl_auto_in_ar_bits_prot),
    .auto_in_r_ready(axi42tl_auto_in_r_ready),
    .auto_in_r_valid(axi42tl_auto_in_r_valid),
    .auto_in_r_bits_id(axi42tl_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi42tl_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi42tl_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi42tl_auto_in_r_bits_last),
    .auto_out_a_ready(axi42tl_auto_out_a_ready),
    .auto_out_a_valid(axi42tl_auto_out_a_valid),
    .auto_out_a_bits_opcode(axi42tl_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(axi42tl_auto_out_a_bits_size),
    .auto_out_a_bits_source(axi42tl_auto_out_a_bits_source),
    .auto_out_a_bits_address(axi42tl_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(axi42tl_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(axi42tl_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(axi42tl_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(axi42tl_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(axi42tl_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(axi42tl_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(axi42tl_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(axi42tl_auto_out_a_bits_mask),
    .auto_out_a_bits_data(axi42tl_auto_out_a_bits_data),
    .auto_out_d_ready(axi42tl_auto_out_d_ready),
    .auto_out_d_valid(axi42tl_auto_out_d_valid),
    .auto_out_d_bits_opcode(axi42tl_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(axi42tl_auto_out_d_bits_size),
    .auto_out_d_bits_source(axi42tl_auto_out_d_bits_source),
    .auto_out_d_bits_denied(axi42tl_auto_out_d_bits_denied),
    .auto_out_d_bits_data(axi42tl_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(axi42tl_auto_out_d_bits_corrupt),
    .io_covSum(axi42tl_io_covSum),
    .metaReset(axi42tl_metaReset)
  );
  AXI4UserYanker axi4yank ( // @[UserYanker.scala 105:30]
    .clock(axi4yank_clock),
    .reset(axi4yank_reset),
    .auto_in_aw_ready(axi4yank_auto_in_aw_ready),
    .auto_in_aw_valid(axi4yank_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4yank_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4yank_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4yank_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4yank_auto_in_aw_bits_size),
    .auto_in_aw_bits_cache(axi4yank_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4yank_auto_in_aw_bits_prot),
    .auto_in_aw_bits_echo_extra_id(axi4yank_auto_in_aw_bits_echo_extra_id),
    .auto_in_aw_bits_echo_real_last(axi4yank_auto_in_aw_bits_echo_real_last),
    .auto_in_w_ready(axi4yank_auto_in_w_ready),
    .auto_in_w_valid(axi4yank_auto_in_w_valid),
    .auto_in_w_bits_data(axi4yank_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4yank_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4yank_auto_in_w_bits_last),
    .auto_in_b_ready(axi4yank_auto_in_b_ready),
    .auto_in_b_valid(axi4yank_auto_in_b_valid),
    .auto_in_b_bits_id(axi4yank_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4yank_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_extra_id(axi4yank_auto_in_b_bits_echo_extra_id),
    .auto_in_b_bits_echo_real_last(axi4yank_auto_in_b_bits_echo_real_last),
    .auto_in_ar_ready(axi4yank_auto_in_ar_ready),
    .auto_in_ar_valid(axi4yank_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4yank_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4yank_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4yank_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4yank_auto_in_ar_bits_size),
    .auto_in_ar_bits_cache(axi4yank_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4yank_auto_in_ar_bits_prot),
    .auto_in_ar_bits_echo_extra_id(axi4yank_auto_in_ar_bits_echo_extra_id),
    .auto_in_ar_bits_echo_real_last(axi4yank_auto_in_ar_bits_echo_real_last),
    .auto_in_r_ready(axi4yank_auto_in_r_ready),
    .auto_in_r_valid(axi4yank_auto_in_r_valid),
    .auto_in_r_bits_id(axi4yank_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4yank_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4yank_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_extra_id(axi4yank_auto_in_r_bits_echo_extra_id),
    .auto_in_r_bits_echo_real_last(axi4yank_auto_in_r_bits_echo_real_last),
    .auto_in_r_bits_last(axi4yank_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4yank_auto_out_aw_ready),
    .auto_out_aw_valid(axi4yank_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4yank_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4yank_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4yank_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4yank_auto_out_aw_bits_size),
    .auto_out_aw_bits_cache(axi4yank_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4yank_auto_out_aw_bits_prot),
    .auto_out_w_ready(axi4yank_auto_out_w_ready),
    .auto_out_w_valid(axi4yank_auto_out_w_valid),
    .auto_out_w_bits_data(axi4yank_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4yank_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4yank_auto_out_w_bits_last),
    .auto_out_b_ready(axi4yank_auto_out_b_ready),
    .auto_out_b_valid(axi4yank_auto_out_b_valid),
    .auto_out_b_bits_id(axi4yank_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4yank_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4yank_auto_out_ar_ready),
    .auto_out_ar_valid(axi4yank_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4yank_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4yank_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4yank_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4yank_auto_out_ar_bits_size),
    .auto_out_ar_bits_cache(axi4yank_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4yank_auto_out_ar_bits_prot),
    .auto_out_r_ready(axi4yank_auto_out_r_ready),
    .auto_out_r_valid(axi4yank_auto_out_r_valid),
    .auto_out_r_bits_id(axi4yank_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4yank_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4yank_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4yank_auto_out_r_bits_last),
    .io_covSum(axi4yank_io_covSum)
  );
  AXI4Fragmenter axi4frag ( // @[Fragmenter.scala 205:30]
    .clock(axi4frag_clock),
    .reset(axi4frag_reset),
    .auto_in_aw_ready(axi4frag_auto_in_aw_ready),
    .auto_in_aw_valid(axi4frag_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4frag_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4frag_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4frag_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4frag_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4frag_auto_in_aw_bits_burst),
    .auto_in_aw_bits_cache(axi4frag_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4frag_auto_in_aw_bits_prot),
    .auto_in_aw_bits_echo_extra_id(axi4frag_auto_in_aw_bits_echo_extra_id),
    .auto_in_w_ready(axi4frag_auto_in_w_ready),
    .auto_in_w_valid(axi4frag_auto_in_w_valid),
    .auto_in_w_bits_data(axi4frag_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4frag_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4frag_auto_in_w_bits_last),
    .auto_in_b_ready(axi4frag_auto_in_b_ready),
    .auto_in_b_valid(axi4frag_auto_in_b_valid),
    .auto_in_b_bits_id(axi4frag_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4frag_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_extra_id(axi4frag_auto_in_b_bits_echo_extra_id),
    .auto_in_ar_ready(axi4frag_auto_in_ar_ready),
    .auto_in_ar_valid(axi4frag_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4frag_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4frag_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4frag_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4frag_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4frag_auto_in_ar_bits_burst),
    .auto_in_ar_bits_cache(axi4frag_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4frag_auto_in_ar_bits_prot),
    .auto_in_ar_bits_echo_extra_id(axi4frag_auto_in_ar_bits_echo_extra_id),
    .auto_in_r_ready(axi4frag_auto_in_r_ready),
    .auto_in_r_valid(axi4frag_auto_in_r_valid),
    .auto_in_r_bits_id(axi4frag_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4frag_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4frag_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_extra_id(axi4frag_auto_in_r_bits_echo_extra_id),
    .auto_in_r_bits_last(axi4frag_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4frag_auto_out_aw_ready),
    .auto_out_aw_valid(axi4frag_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4frag_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4frag_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4frag_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4frag_auto_out_aw_bits_size),
    .auto_out_aw_bits_cache(axi4frag_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4frag_auto_out_aw_bits_prot),
    .auto_out_aw_bits_echo_extra_id(axi4frag_auto_out_aw_bits_echo_extra_id),
    .auto_out_aw_bits_echo_real_last(axi4frag_auto_out_aw_bits_echo_real_last),
    .auto_out_w_ready(axi4frag_auto_out_w_ready),
    .auto_out_w_valid(axi4frag_auto_out_w_valid),
    .auto_out_w_bits_data(axi4frag_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4frag_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4frag_auto_out_w_bits_last),
    .auto_out_b_ready(axi4frag_auto_out_b_ready),
    .auto_out_b_valid(axi4frag_auto_out_b_valid),
    .auto_out_b_bits_id(axi4frag_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4frag_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_extra_id(axi4frag_auto_out_b_bits_echo_extra_id),
    .auto_out_b_bits_echo_real_last(axi4frag_auto_out_b_bits_echo_real_last),
    .auto_out_ar_ready(axi4frag_auto_out_ar_ready),
    .auto_out_ar_valid(axi4frag_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4frag_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4frag_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4frag_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4frag_auto_out_ar_bits_size),
    .auto_out_ar_bits_cache(axi4frag_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4frag_auto_out_ar_bits_prot),
    .auto_out_ar_bits_echo_extra_id(axi4frag_auto_out_ar_bits_echo_extra_id),
    .auto_out_ar_bits_echo_real_last(axi4frag_auto_out_ar_bits_echo_real_last),
    .auto_out_r_ready(axi4frag_auto_out_r_ready),
    .auto_out_r_valid(axi4frag_auto_out_r_valid),
    .auto_out_r_bits_id(axi4frag_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4frag_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4frag_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_extra_id(axi4frag_auto_out_r_bits_echo_extra_id),
    .auto_out_r_bits_echo_real_last(axi4frag_auto_out_r_bits_echo_real_last),
    .auto_out_r_bits_last(axi4frag_auto_out_r_bits_last),
    .io_covSum(axi4frag_io_covSum),
    .metaReset(axi4frag_metaReset)
  );
  AXI4IdIndexer axi4index ( // @[IdIndexer.scala 91:31]
    .auto_in_aw_ready(axi4index_auto_in_aw_ready),
    .auto_in_aw_valid(axi4index_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4index_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4index_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4index_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4index_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4index_auto_in_aw_bits_burst),
    .auto_in_aw_bits_cache(axi4index_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4index_auto_in_aw_bits_prot),
    .auto_in_w_ready(axi4index_auto_in_w_ready),
    .auto_in_w_valid(axi4index_auto_in_w_valid),
    .auto_in_w_bits_data(axi4index_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4index_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4index_auto_in_w_bits_last),
    .auto_in_b_ready(axi4index_auto_in_b_ready),
    .auto_in_b_valid(axi4index_auto_in_b_valid),
    .auto_in_b_bits_id(axi4index_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4index_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4index_auto_in_ar_ready),
    .auto_in_ar_valid(axi4index_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4index_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4index_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4index_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4index_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4index_auto_in_ar_bits_burst),
    .auto_in_ar_bits_cache(axi4index_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4index_auto_in_ar_bits_prot),
    .auto_in_r_ready(axi4index_auto_in_r_ready),
    .auto_in_r_valid(axi4index_auto_in_r_valid),
    .auto_in_r_bits_id(axi4index_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4index_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4index_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4index_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4index_auto_out_aw_ready),
    .auto_out_aw_valid(axi4index_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4index_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4index_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4index_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4index_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4index_auto_out_aw_bits_burst),
    .auto_out_aw_bits_cache(axi4index_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4index_auto_out_aw_bits_prot),
    .auto_out_aw_bits_echo_extra_id(axi4index_auto_out_aw_bits_echo_extra_id),
    .auto_out_w_ready(axi4index_auto_out_w_ready),
    .auto_out_w_valid(axi4index_auto_out_w_valid),
    .auto_out_w_bits_data(axi4index_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4index_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4index_auto_out_w_bits_last),
    .auto_out_b_ready(axi4index_auto_out_b_ready),
    .auto_out_b_valid(axi4index_auto_out_b_valid),
    .auto_out_b_bits_id(axi4index_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4index_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_extra_id(axi4index_auto_out_b_bits_echo_extra_id),
    .auto_out_ar_ready(axi4index_auto_out_ar_ready),
    .auto_out_ar_valid(axi4index_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4index_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4index_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4index_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4index_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4index_auto_out_ar_bits_burst),
    .auto_out_ar_bits_cache(axi4index_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4index_auto_out_ar_bits_prot),
    .auto_out_ar_bits_echo_extra_id(axi4index_auto_out_ar_bits_echo_extra_id),
    .auto_out_r_ready(axi4index_auto_out_r_ready),
    .auto_out_r_valid(axi4index_auto_out_r_valid),
    .auto_out_r_bits_id(axi4index_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4index_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4index_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_extra_id(axi4index_auto_out_r_bits_echo_extra_id),
    .auto_out_r_bits_last(axi4index_auto_out_r_bits_last),
    .io_covSum(axi4index_io_covSum)
  );
  assign widget_auto_in_a_ready = widget_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_valid = widget_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_opcode = widget_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_size = widget_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_source = widget_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_denied = widget_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_data = widget_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_corrupt = widget_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_out_a_valid = widget_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_opcode = widget_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_size = widget_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_source = widget_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_address = widget_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_bufferable = widget_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_modifiable = widget_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_readalloc = widget_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_writealloc = widget_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_privileged = widget_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_secure = widget_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_fetch = widget_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_mask = widget_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_data = widget_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_d_ready = widget_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_axi4index_in_aw_ready = axi4index_auto_in_aw_ready; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_w_ready = axi4index_auto_in_w_ready; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_b_valid = axi4index_auto_in_b_valid; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_b_bits_id = axi4index_auto_in_b_bits_id; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_b_bits_resp = axi4index_auto_in_b_bits_resp; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_ar_ready = axi4index_auto_in_ar_ready; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_r_valid = axi4index_auto_in_r_valid; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_r_bits_id = axi4index_auto_in_r_bits_id; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_r_bits_data = axi4index_auto_in_r_bits_data; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_r_bits_resp = axi4index_auto_in_r_bits_resp; // @[LazyModule.scala 309:16]
  assign auto_axi4index_in_r_bits_last = axi4index_auto_in_r_bits_last; // @[LazyModule.scala 309:16]
  assign auto_tl_out_a_valid = buffer_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_param = buffer_auto_out_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_size = buffer_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_source = buffer_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_address = buffer_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_user_amba_prot_bufferable = buffer_auto_out_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_user_amba_prot_modifiable = buffer_auto_out_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_user_amba_prot_readalloc = buffer_auto_out_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_user_amba_prot_writealloc = buffer_auto_out_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_user_amba_prot_privileged = buffer_auto_out_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_user_amba_prot_secure = buffer_auto_out_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_user_amba_prot_fetch = buffer_auto_out_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_mask = buffer_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_a_bits_data = buffer_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_out_d_ready = buffer_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_a_valid = fixer_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_param = 3'h0; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_size = fixer_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_source = fixer_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_address = fixer_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_bufferable = fixer_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_modifiable = fixer_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_readalloc = fixer_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_writealloc = fixer_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_privileged = fixer_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_secure = fixer_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_fetch = fixer_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_data = fixer_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_d_ready = fixer_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_a_ready = auto_tl_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_d_valid = auto_tl_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_d_bits_opcode = auto_tl_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_d_bits_size = auto_tl_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_d_bits_source = auto_tl_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_d_bits_denied = auto_tl_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_d_bits_data = auto_tl_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_d_bits_corrupt = auto_tl_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign fixer_clock = clock;
  assign fixer_reset = reset;
  assign fixer_auto_in_a_valid = widget_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_size = widget_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_source = widget_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_address = widget_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_bufferable = widget_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_modifiable = widget_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_readalloc = widget_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_writealloc = widget_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_privileged = widget_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_secure = widget_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_fetch = widget_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_mask = widget_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_data = widget_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_d_ready = widget_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_valid = axi42tl_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_opcode = axi42tl_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_size = axi42tl_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_source = axi42tl_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_address = axi42tl_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_bufferable = axi42tl_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_modifiable = axi42tl_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_readalloc = axi42tl_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_writealloc = axi42tl_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_privileged = axi42tl_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_secure = axi42tl_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_fetch = axi42tl_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_mask = axi42tl_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_data = axi42tl_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign widget_auto_in_d_ready = axi42tl_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign widget_auto_out_a_ready = fixer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_valid = fixer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_size = fixer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_source = fixer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_denied = fixer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_data = fixer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign axi42tl_clock = clock;
  assign axi42tl_reset = reset;
  assign axi42tl_auto_in_aw_valid = axi4yank_auto_out_aw_valid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_id = axi4yank_auto_out_aw_bits_id; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_addr = axi4yank_auto_out_aw_bits_addr; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_len = axi4yank_auto_out_aw_bits_len; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_size = axi4yank_auto_out_aw_bits_size; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_cache = axi4yank_auto_out_aw_bits_cache; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_prot = axi4yank_auto_out_aw_bits_prot; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_w_valid = axi4yank_auto_out_w_valid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_w_bits_data = axi4yank_auto_out_w_bits_data; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_w_bits_strb = axi4yank_auto_out_w_bits_strb; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_w_bits_last = axi4yank_auto_out_w_bits_last; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_b_ready = axi4yank_auto_out_b_ready; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_valid = axi4yank_auto_out_ar_valid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_id = axi4yank_auto_out_ar_bits_id; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_addr = axi4yank_auto_out_ar_bits_addr; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_len = axi4yank_auto_out_ar_bits_len; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_size = axi4yank_auto_out_ar_bits_size; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_cache = axi4yank_auto_out_ar_bits_cache; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_prot = axi4yank_auto_out_ar_bits_prot; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_r_ready = axi4yank_auto_out_r_ready; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_a_ready = widget_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_valid = widget_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_opcode = widget_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_size = widget_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_source = widget_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_denied = widget_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_data = widget_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_corrupt = widget_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign axi4yank_clock = clock;
  assign axi4yank_reset = reset;
  assign axi4yank_auto_in_aw_valid = axi4frag_auto_out_aw_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_id = axi4frag_auto_out_aw_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_addr = axi4frag_auto_out_aw_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_len = axi4frag_auto_out_aw_bits_len; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_size = axi4frag_auto_out_aw_bits_size; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_cache = axi4frag_auto_out_aw_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_prot = axi4frag_auto_out_aw_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_echo_extra_id = axi4frag_auto_out_aw_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_echo_real_last = axi4frag_auto_out_aw_bits_echo_real_last; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_valid = axi4frag_auto_out_w_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_bits_data = axi4frag_auto_out_w_bits_data; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_bits_strb = axi4frag_auto_out_w_bits_strb; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_bits_last = axi4frag_auto_out_w_bits_last; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_b_ready = axi4frag_auto_out_b_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_valid = axi4frag_auto_out_ar_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_id = axi4frag_auto_out_ar_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_addr = axi4frag_auto_out_ar_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_len = axi4frag_auto_out_ar_bits_len; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_size = axi4frag_auto_out_ar_bits_size; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_cache = axi4frag_auto_out_ar_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_prot = axi4frag_auto_out_ar_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_echo_extra_id = axi4frag_auto_out_ar_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_echo_real_last = axi4frag_auto_out_ar_bits_echo_real_last; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_r_ready = axi4frag_auto_out_r_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_aw_ready = axi42tl_auto_in_aw_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_w_ready = axi42tl_auto_in_w_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_b_valid = axi42tl_auto_in_b_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_b_bits_id = axi42tl_auto_in_b_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_b_bits_resp = axi42tl_auto_in_b_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_ar_ready = axi42tl_auto_in_ar_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_valid = axi42tl_auto_in_r_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_bits_id = axi42tl_auto_in_r_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_bits_data = axi42tl_auto_in_r_bits_data; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_bits_resp = axi42tl_auto_in_r_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_bits_last = axi42tl_auto_in_r_bits_last; // @[LazyModule.scala 296:16]
  assign axi4frag_clock = clock;
  assign axi4frag_reset = reset;
  assign axi4frag_auto_in_aw_valid = axi4index_auto_out_aw_valid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_aw_bits_id = axi4index_auto_out_aw_bits_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_aw_bits_addr = axi4index_auto_out_aw_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_aw_bits_len = axi4index_auto_out_aw_bits_len; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_aw_bits_size = axi4index_auto_out_aw_bits_size; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_aw_bits_burst = axi4index_auto_out_aw_bits_burst; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_aw_bits_cache = axi4index_auto_out_aw_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_aw_bits_prot = axi4index_auto_out_aw_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_aw_bits_echo_extra_id = axi4index_auto_out_aw_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_w_valid = axi4index_auto_out_w_valid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_w_bits_data = axi4index_auto_out_w_bits_data; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_w_bits_strb = axi4index_auto_out_w_bits_strb; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_w_bits_last = axi4index_auto_out_w_bits_last; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_b_ready = axi4index_auto_out_b_ready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_ar_valid = axi4index_auto_out_ar_valid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_ar_bits_id = axi4index_auto_out_ar_bits_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_ar_bits_addr = axi4index_auto_out_ar_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_ar_bits_len = axi4index_auto_out_ar_bits_len; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_ar_bits_size = axi4index_auto_out_ar_bits_size; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_ar_bits_burst = axi4index_auto_out_ar_bits_burst; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_ar_bits_cache = axi4index_auto_out_ar_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_ar_bits_prot = axi4index_auto_out_ar_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_ar_bits_echo_extra_id = axi4index_auto_out_ar_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_in_r_ready = axi4index_auto_out_r_ready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_aw_ready = axi4yank_auto_in_aw_ready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_w_ready = axi4yank_auto_in_w_ready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_b_valid = axi4yank_auto_in_b_valid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_b_bits_id = axi4yank_auto_in_b_bits_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_b_bits_resp = axi4yank_auto_in_b_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_b_bits_echo_extra_id = axi4yank_auto_in_b_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_b_bits_echo_real_last = axi4yank_auto_in_b_bits_echo_real_last; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_ar_ready = axi4yank_auto_in_ar_ready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_valid = axi4yank_auto_in_r_valid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_id = axi4yank_auto_in_r_bits_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_data = axi4yank_auto_in_r_bits_data; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_resp = axi4yank_auto_in_r_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_echo_extra_id = axi4yank_auto_in_r_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_echo_real_last = axi4yank_auto_in_r_bits_echo_real_last; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_last = axi4yank_auto_in_r_bits_last; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_valid = auto_axi4index_in_aw_valid; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_aw_bits_id = auto_axi4index_in_aw_bits_id; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_aw_bits_addr = auto_axi4index_in_aw_bits_addr; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_aw_bits_len = auto_axi4index_in_aw_bits_len; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_aw_bits_size = auto_axi4index_in_aw_bits_size; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_aw_bits_burst = auto_axi4index_in_aw_bits_burst; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_aw_bits_cache = auto_axi4index_in_aw_bits_cache; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_aw_bits_prot = auto_axi4index_in_aw_bits_prot; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_w_valid = auto_axi4index_in_w_valid; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_w_bits_data = auto_axi4index_in_w_bits_data; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_w_bits_strb = auto_axi4index_in_w_bits_strb; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_w_bits_last = auto_axi4index_in_w_bits_last; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_b_ready = auto_axi4index_in_b_ready; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_ar_valid = auto_axi4index_in_ar_valid; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_ar_bits_id = auto_axi4index_in_ar_bits_id; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_ar_bits_addr = auto_axi4index_in_ar_bits_addr; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_ar_bits_len = auto_axi4index_in_ar_bits_len; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_ar_bits_size = auto_axi4index_in_ar_bits_size; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_ar_bits_burst = auto_axi4index_in_ar_bits_burst; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_ar_bits_cache = auto_axi4index_in_ar_bits_cache; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_ar_bits_prot = auto_axi4index_in_ar_bits_prot; // @[LazyModule.scala 309:16]
  assign axi4index_auto_in_r_ready = auto_axi4index_in_r_ready; // @[LazyModule.scala 309:16]
  assign axi4index_auto_out_aw_ready = axi4frag_auto_in_aw_ready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_w_ready = axi4frag_auto_in_w_ready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_valid = axi4frag_auto_in_b_valid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_bits_id = axi4frag_auto_in_b_bits_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_bits_resp = axi4frag_auto_in_b_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_bits_echo_extra_id = axi4frag_auto_in_b_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_ar_ready = axi4frag_auto_in_ar_ready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_valid = axi4frag_auto_in_r_valid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_id = axi4frag_auto_in_r_bits_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_data = axi4frag_auto_in_r_bits_data; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_resp = axi4frag_auto_in_r_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_echo_extra_id = axi4frag_auto_in_r_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_last = axi4frag_auto_in_r_bits_last; // @[LazyModule.scala 296:16]
  assign TLInterconnectCoupler_5_covSum = 30'h0;
  assign fixer_sum = TLInterconnectCoupler_5_covSum + fixer_io_covSum;
  assign axi42tl_sum = fixer_sum + axi42tl_io_covSum;
  assign axi4yank_sum = axi42tl_sum + axi4yank_io_covSum;
  assign axi4frag_sum = axi4yank_sum + axi4frag_io_covSum;
  assign buffer_sum = axi4frag_sum + buffer_io_covSum;
  assign axi4index_sum = buffer_sum + axi4index_io_covSum;
  assign io_covSum = axi4index_sum;
  assign fixer_metaReset = metaReset;
  assign axi42tl_metaReset = metaReset;
  assign axi4frag_metaReset = metaReset;
endmodule
module TLFIFOFixer_3(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [30:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [30:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_101;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_102;
`endif // RANDOMIZE_REG_INIT
  wire [30:0] _a_id_T = auto_in_a_bits_address ^ 31'h2000; // @[Parameters.scala 137:31]
  wire [31:0] _a_id_T_1 = {1'b0,$signed(_a_id_T)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_id_T_3 = $signed(_a_id_T_1) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  _a_id_T_4 = $signed(_a_id_T_3) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _a_id_T_5 = auto_in_a_bits_address ^ 31'h44000000; // @[Parameters.scala 137:31]
  wire [31:0] _a_id_T_6 = {1'b0,$signed(_a_id_T_5)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_id_T_8 = $signed(_a_id_T_6) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  _a_id_T_9 = $signed(_a_id_T_8) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _a_id_T_10 = auto_in_a_bits_address ^ 31'h4000000; // @[Parameters.scala 137:31]
  wire [31:0] _a_id_T_11 = {1'b0,$signed(_a_id_T_10)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_id_T_13 = $signed(_a_id_T_11) & 32'sh44000000; // @[Parameters.scala 137:52]
  wire  _a_id_T_14 = $signed(_a_id_T_13) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _a_id_T_15 = auto_in_a_bits_address ^ 31'h2000000; // @[Parameters.scala 137:31]
  wire [31:0] _a_id_T_16 = {1'b0,$signed(_a_id_T_15)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_id_T_18 = $signed(_a_id_T_16) & 32'sh46030000; // @[Parameters.scala 137:52]
  wire  _a_id_T_19 = $signed(_a_id_T_18) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _a_id_T_20 = auto_in_a_bits_address ^ 31'h10000; // @[Parameters.scala 137:31]
  wire [31:0] _a_id_T_21 = {1'b0,$signed(_a_id_T_20)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_id_T_23 = $signed(_a_id_T_21) & 32'sh46030000; // @[Parameters.scala 137:52]
  wire  _a_id_T_24 = $signed(_a_id_T_23) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _a_id_T_25 = auto_in_a_bits_address ^ 31'h20000; // @[Parameters.scala 137:31]
  wire [31:0] _a_id_T_26 = {1'b0,$signed(_a_id_T_25)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_id_T_28 = $signed(_a_id_T_26) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  _a_id_T_29 = $signed(_a_id_T_28) == 32'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _a_id_T_31 = {1'b0,$signed(auto_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_id_T_33 = $signed(_a_id_T_31) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  _a_id_T_34 = $signed(_a_id_T_33) == 32'sh0; // @[Parameters.scala 137:67]
  wire [1:0] _a_id_T_36 = _a_id_T_9 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _a_id_T_37 = _a_id_T_14 ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _a_id_T_38 = _a_id_T_19 ? 3'h6 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _a_id_T_39 = _a_id_T_24 ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [1:0] _a_id_T_40 = _a_id_T_29 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _a_id_T_41 = _a_id_T_34 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_340 = {{1'd0}, _a_id_T_4}; // @[Mux.scala 27:73]
  wire [1:0] _a_id_T_42 = _GEN_340 | _a_id_T_36; // @[Mux.scala 27:73]
  wire [2:0] _GEN_341 = {{1'd0}, _a_id_T_42}; // @[Mux.scala 27:73]
  wire [2:0] _a_id_T_43 = _GEN_341 | _a_id_T_37; // @[Mux.scala 27:73]
  wire [2:0] _a_id_T_44 = _a_id_T_43 | _a_id_T_38; // @[Mux.scala 27:73]
  wire [2:0] _a_id_T_45 = _a_id_T_44 | _a_id_T_39; // @[Mux.scala 27:73]
  wire [2:0] _GEN_342 = {{1'd0}, _a_id_T_40}; // @[Mux.scala 27:73]
  wire [2:0] _a_id_T_46 = _a_id_T_45 | _GEN_342; // @[Mux.scala 27:73]
  wire [2:0] a_id = _a_id_T_46 | _a_id_T_41; // @[Mux.scala 27:73]
  wire  a_noDomain = a_id == 3'h0; // @[FIFOFixer.scala 55:29]
  wire  stalls_a_sel = auto_in_a_bits_source[6:3] == 4'h8; // @[Parameters.scala 54:32]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25]
  reg  flight_64; // @[FIFOFixer.scala 71:27]
  reg  flight_65; // @[FIFOFixer.scala 71:27]
  reg  flight_66; // @[FIFOFixer.scala 71:27]
  reg  flight_67; // @[FIFOFixer.scala 71:27]
  reg  flight_68; // @[FIFOFixer.scala 71:27]
  reg  flight_69; // @[FIFOFixer.scala 71:27]
  reg  flight_70; // @[FIFOFixer.scala 71:27]
  reg  flight_71; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id; // @[Reg.scala 16:16]
  wire  stalls_0 = stalls_a_sel & a_first & (flight_64 | flight_65 | flight_66 | flight_67 | flight_68 | flight_69 |
    flight_70 | flight_71) & (a_noDomain | stalls_id != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_1 = auto_in_a_bits_source[6:3] == 4'h9; // @[Parameters.scala 54:32]
  reg  flight_72; // @[FIFOFixer.scala 71:27]
  reg  flight_73; // @[FIFOFixer.scala 71:27]
  reg  flight_74; // @[FIFOFixer.scala 71:27]
  reg  flight_75; // @[FIFOFixer.scala 71:27]
  reg  flight_76; // @[FIFOFixer.scala 71:27]
  reg  flight_77; // @[FIFOFixer.scala 71:27]
  reg  flight_78; // @[FIFOFixer.scala 71:27]
  reg  flight_79; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_1; // @[Reg.scala 16:16]
  wire  stalls_1 = stalls_a_sel_1 & a_first & (flight_72 | flight_73 | flight_74 | flight_75 | flight_76 | flight_77 |
    flight_78 | flight_79) & (a_noDomain | stalls_id_1 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_2 = auto_in_a_bits_source[6:2] == 5'h0; // @[Parameters.scala 54:32]
  reg  flight_0; // @[FIFOFixer.scala 71:27]
  reg  flight_1; // @[FIFOFixer.scala 71:27]
  reg  flight_2; // @[FIFOFixer.scala 71:27]
  reg  flight_3; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_2; // @[Reg.scala 16:16]
  wire  stalls_2 = stalls_a_sel_2 & a_first & (flight_0 | flight_1 | flight_2 | flight_3) & (a_noDomain | stalls_id_2
     != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_3 = auto_in_a_bits_source[6:2] == 5'h1; // @[Parameters.scala 54:32]
  reg  flight_4; // @[FIFOFixer.scala 71:27]
  reg  flight_5; // @[FIFOFixer.scala 71:27]
  reg  flight_6; // @[FIFOFixer.scala 71:27]
  reg  flight_7; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_3; // @[Reg.scala 16:16]
  wire  stalls_3 = stalls_a_sel_3 & a_first & (flight_4 | flight_5 | flight_6 | flight_7) & (a_noDomain | stalls_id_3
     != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_4 = auto_in_a_bits_source[6:2] == 5'h2; // @[Parameters.scala 54:32]
  reg  flight_8; // @[FIFOFixer.scala 71:27]
  reg  flight_9; // @[FIFOFixer.scala 71:27]
  reg  flight_10; // @[FIFOFixer.scala 71:27]
  reg  flight_11; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_4; // @[Reg.scala 16:16]
  wire  stalls_4 = stalls_a_sel_4 & a_first & (flight_8 | flight_9 | flight_10 | flight_11) & (a_noDomain | stalls_id_4
     != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_5 = auto_in_a_bits_source[6:2] == 5'h3; // @[Parameters.scala 54:32]
  reg  flight_12; // @[FIFOFixer.scala 71:27]
  reg  flight_13; // @[FIFOFixer.scala 71:27]
  reg  flight_14; // @[FIFOFixer.scala 71:27]
  reg  flight_15; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_5; // @[Reg.scala 16:16]
  wire  stalls_5 = stalls_a_sel_5 & a_first & (flight_12 | flight_13 | flight_14 | flight_15) & (a_noDomain |
    stalls_id_5 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_6 = auto_in_a_bits_source[6:2] == 5'h4; // @[Parameters.scala 54:32]
  reg  flight_16; // @[FIFOFixer.scala 71:27]
  reg  flight_17; // @[FIFOFixer.scala 71:27]
  reg  flight_18; // @[FIFOFixer.scala 71:27]
  reg  flight_19; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_6; // @[Reg.scala 16:16]
  wire  stalls_6 = stalls_a_sel_6 & a_first & (flight_16 | flight_17 | flight_18 | flight_19) & (a_noDomain |
    stalls_id_6 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_7 = auto_in_a_bits_source[6:2] == 5'h5; // @[Parameters.scala 54:32]
  reg  flight_20; // @[FIFOFixer.scala 71:27]
  reg  flight_21; // @[FIFOFixer.scala 71:27]
  reg  flight_22; // @[FIFOFixer.scala 71:27]
  reg  flight_23; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_7; // @[Reg.scala 16:16]
  wire  stalls_7 = stalls_a_sel_7 & a_first & (flight_20 | flight_21 | flight_22 | flight_23) & (a_noDomain |
    stalls_id_7 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_8 = auto_in_a_bits_source[6:2] == 5'h6; // @[Parameters.scala 54:32]
  reg  flight_24; // @[FIFOFixer.scala 71:27]
  reg  flight_25; // @[FIFOFixer.scala 71:27]
  reg  flight_26; // @[FIFOFixer.scala 71:27]
  reg  flight_27; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_8; // @[Reg.scala 16:16]
  wire  stalls_8 = stalls_a_sel_8 & a_first & (flight_24 | flight_25 | flight_26 | flight_27) & (a_noDomain |
    stalls_id_8 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_9 = auto_in_a_bits_source[6:2] == 5'h7; // @[Parameters.scala 54:32]
  reg  flight_28; // @[FIFOFixer.scala 71:27]
  reg  flight_29; // @[FIFOFixer.scala 71:27]
  reg  flight_30; // @[FIFOFixer.scala 71:27]
  reg  flight_31; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_9; // @[Reg.scala 16:16]
  wire  stalls_9 = stalls_a_sel_9 & a_first & (flight_28 | flight_29 | flight_30 | flight_31) & (a_noDomain |
    stalls_id_9 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_10 = auto_in_a_bits_source[6:2] == 5'h8; // @[Parameters.scala 54:32]
  reg  flight_32; // @[FIFOFixer.scala 71:27]
  reg  flight_33; // @[FIFOFixer.scala 71:27]
  reg  flight_34; // @[FIFOFixer.scala 71:27]
  reg  flight_35; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_10; // @[Reg.scala 16:16]
  wire  stalls_10 = stalls_a_sel_10 & a_first & (flight_32 | flight_33 | flight_34 | flight_35) & (a_noDomain |
    stalls_id_10 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_11 = auto_in_a_bits_source[6:2] == 5'h9; // @[Parameters.scala 54:32]
  reg  flight_36; // @[FIFOFixer.scala 71:27]
  reg  flight_37; // @[FIFOFixer.scala 71:27]
  reg  flight_38; // @[FIFOFixer.scala 71:27]
  reg  flight_39; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_11; // @[Reg.scala 16:16]
  wire  stalls_11 = stalls_a_sel_11 & a_first & (flight_36 | flight_37 | flight_38 | flight_39) & (a_noDomain |
    stalls_id_11 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_12 = auto_in_a_bits_source[6:2] == 5'ha; // @[Parameters.scala 54:32]
  reg  flight_40; // @[FIFOFixer.scala 71:27]
  reg  flight_41; // @[FIFOFixer.scala 71:27]
  reg  flight_42; // @[FIFOFixer.scala 71:27]
  reg  flight_43; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_12; // @[Reg.scala 16:16]
  wire  stalls_12 = stalls_a_sel_12 & a_first & (flight_40 | flight_41 | flight_42 | flight_43) & (a_noDomain |
    stalls_id_12 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_13 = auto_in_a_bits_source[6:2] == 5'hb; // @[Parameters.scala 54:32]
  reg  flight_44; // @[FIFOFixer.scala 71:27]
  reg  flight_45; // @[FIFOFixer.scala 71:27]
  reg  flight_46; // @[FIFOFixer.scala 71:27]
  reg  flight_47; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_13; // @[Reg.scala 16:16]
  wire  stalls_13 = stalls_a_sel_13 & a_first & (flight_44 | flight_45 | flight_46 | flight_47) & (a_noDomain |
    stalls_id_13 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_14 = auto_in_a_bits_source[6:2] == 5'hc; // @[Parameters.scala 54:32]
  reg  flight_48; // @[FIFOFixer.scala 71:27]
  reg  flight_49; // @[FIFOFixer.scala 71:27]
  reg  flight_50; // @[FIFOFixer.scala 71:27]
  reg  flight_51; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_14; // @[Reg.scala 16:16]
  wire  stalls_14 = stalls_a_sel_14 & a_first & (flight_48 | flight_49 | flight_50 | flight_51) & (a_noDomain |
    stalls_id_14 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_15 = auto_in_a_bits_source[6:2] == 5'hd; // @[Parameters.scala 54:32]
  reg  flight_52; // @[FIFOFixer.scala 71:27]
  reg  flight_53; // @[FIFOFixer.scala 71:27]
  reg  flight_54; // @[FIFOFixer.scala 71:27]
  reg  flight_55; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_15; // @[Reg.scala 16:16]
  wire  stalls_15 = stalls_a_sel_15 & a_first & (flight_52 | flight_53 | flight_54 | flight_55) & (a_noDomain |
    stalls_id_15 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_16 = auto_in_a_bits_source[6:2] == 5'he; // @[Parameters.scala 54:32]
  reg  flight_56; // @[FIFOFixer.scala 71:27]
  reg  flight_57; // @[FIFOFixer.scala 71:27]
  reg  flight_58; // @[FIFOFixer.scala 71:27]
  reg  flight_59; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_16; // @[Reg.scala 16:16]
  wire  stalls_16 = stalls_a_sel_16 & a_first & (flight_56 | flight_57 | flight_58 | flight_59) & (a_noDomain |
    stalls_id_16 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_17 = auto_in_a_bits_source[6:2] == 5'hf; // @[Parameters.scala 54:32]
  reg  flight_60; // @[FIFOFixer.scala 71:27]
  reg  flight_61; // @[FIFOFixer.scala 71:27]
  reg  flight_62; // @[FIFOFixer.scala 71:27]
  reg  flight_63; // @[FIFOFixer.scala 71:27]
  reg [2:0] stalls_id_17; // @[Reg.scala 16:16]
  wire  stalls_17 = stalls_a_sel_17 & a_first & (flight_60 | flight_61 | flight_62 | flight_63) & (a_noDomain |
    stalls_id_17 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stall = stalls_0 | stalls_1 | stalls_2 | stalls_3 | stalls_4 | stalls_5 | stalls_6 | stalls_7 | stalls_8 |
    stalls_9 | stalls_10 | stalls_11 | stalls_12 | stalls_13 | stalls_14 | stalls_15 | stalls_16 | stalls_17; // @[FIFOFixer.scala 83:49]
  wire  _bundleIn_0_a_ready_T = ~stall; // @[FIFOFixer.scala 88:50]
  wire  bundleIn_0_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  wire  _a_first_T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _a_first_beats1_decode_T_1 = 27'hfff << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [11:0] _a_first_beats1_decode_T_3 = ~_a_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] a_first_beats1_decode = _a_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28]
  wire  _d_first_T = auto_in_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28]
  wire  d_first_first = d_first_counter == 9'h0; // @[Edges.scala 230:25]
  wire  d_first = d_first_first & auto_out_d_bits_opcode != 3'h6; // @[FIFOFixer.scala 67:42]
  wire  _GEN_82 = a_first & _a_first_T ? 7'h0 == auto_in_a_bits_source | flight_0 : flight_0; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_83 = a_first & _a_first_T ? 7'h1 == auto_in_a_bits_source | flight_1 : flight_1; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_84 = a_first & _a_first_T ? 7'h2 == auto_in_a_bits_source | flight_2 : flight_2; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_85 = a_first & _a_first_T ? 7'h3 == auto_in_a_bits_source | flight_3 : flight_3; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_86 = a_first & _a_first_T ? 7'h4 == auto_in_a_bits_source | flight_4 : flight_4; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_87 = a_first & _a_first_T ? 7'h5 == auto_in_a_bits_source | flight_5 : flight_5; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_88 = a_first & _a_first_T ? 7'h6 == auto_in_a_bits_source | flight_6 : flight_6; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_89 = a_first & _a_first_T ? 7'h7 == auto_in_a_bits_source | flight_7 : flight_7; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_90 = a_first & _a_first_T ? 7'h8 == auto_in_a_bits_source | flight_8 : flight_8; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_91 = a_first & _a_first_T ? 7'h9 == auto_in_a_bits_source | flight_9 : flight_9; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_92 = a_first & _a_first_T ? 7'ha == auto_in_a_bits_source | flight_10 : flight_10; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_93 = a_first & _a_first_T ? 7'hb == auto_in_a_bits_source | flight_11 : flight_11; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_94 = a_first & _a_first_T ? 7'hc == auto_in_a_bits_source | flight_12 : flight_12; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_95 = a_first & _a_first_T ? 7'hd == auto_in_a_bits_source | flight_13 : flight_13; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_96 = a_first & _a_first_T ? 7'he == auto_in_a_bits_source | flight_14 : flight_14; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_97 = a_first & _a_first_T ? 7'hf == auto_in_a_bits_source | flight_15 : flight_15; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_98 = a_first & _a_first_T ? 7'h10 == auto_in_a_bits_source | flight_16 : flight_16; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_99 = a_first & _a_first_T ? 7'h11 == auto_in_a_bits_source | flight_17 : flight_17; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_100 = a_first & _a_first_T ? 7'h12 == auto_in_a_bits_source | flight_18 : flight_18; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_101 = a_first & _a_first_T ? 7'h13 == auto_in_a_bits_source | flight_19 : flight_19; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_102 = a_first & _a_first_T ? 7'h14 == auto_in_a_bits_source | flight_20 : flight_20; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_103 = a_first & _a_first_T ? 7'h15 == auto_in_a_bits_source | flight_21 : flight_21; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_104 = a_first & _a_first_T ? 7'h16 == auto_in_a_bits_source | flight_22 : flight_22; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_105 = a_first & _a_first_T ? 7'h17 == auto_in_a_bits_source | flight_23 : flight_23; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_106 = a_first & _a_first_T ? 7'h18 == auto_in_a_bits_source | flight_24 : flight_24; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_107 = a_first & _a_first_T ? 7'h19 == auto_in_a_bits_source | flight_25 : flight_25; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_108 = a_first & _a_first_T ? 7'h1a == auto_in_a_bits_source | flight_26 : flight_26; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_109 = a_first & _a_first_T ? 7'h1b == auto_in_a_bits_source | flight_27 : flight_27; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_110 = a_first & _a_first_T ? 7'h1c == auto_in_a_bits_source | flight_28 : flight_28; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_111 = a_first & _a_first_T ? 7'h1d == auto_in_a_bits_source | flight_29 : flight_29; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_112 = a_first & _a_first_T ? 7'h1e == auto_in_a_bits_source | flight_30 : flight_30; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_113 = a_first & _a_first_T ? 7'h1f == auto_in_a_bits_source | flight_31 : flight_31; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_114 = a_first & _a_first_T ? 7'h20 == auto_in_a_bits_source | flight_32 : flight_32; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_115 = a_first & _a_first_T ? 7'h21 == auto_in_a_bits_source | flight_33 : flight_33; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_116 = a_first & _a_first_T ? 7'h22 == auto_in_a_bits_source | flight_34 : flight_34; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_117 = a_first & _a_first_T ? 7'h23 == auto_in_a_bits_source | flight_35 : flight_35; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_118 = a_first & _a_first_T ? 7'h24 == auto_in_a_bits_source | flight_36 : flight_36; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_119 = a_first & _a_first_T ? 7'h25 == auto_in_a_bits_source | flight_37 : flight_37; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_120 = a_first & _a_first_T ? 7'h26 == auto_in_a_bits_source | flight_38 : flight_38; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_121 = a_first & _a_first_T ? 7'h27 == auto_in_a_bits_source | flight_39 : flight_39; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_122 = a_first & _a_first_T ? 7'h28 == auto_in_a_bits_source | flight_40 : flight_40; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_123 = a_first & _a_first_T ? 7'h29 == auto_in_a_bits_source | flight_41 : flight_41; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_124 = a_first & _a_first_T ? 7'h2a == auto_in_a_bits_source | flight_42 : flight_42; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_125 = a_first & _a_first_T ? 7'h2b == auto_in_a_bits_source | flight_43 : flight_43; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_126 = a_first & _a_first_T ? 7'h2c == auto_in_a_bits_source | flight_44 : flight_44; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_127 = a_first & _a_first_T ? 7'h2d == auto_in_a_bits_source | flight_45 : flight_45; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_128 = a_first & _a_first_T ? 7'h2e == auto_in_a_bits_source | flight_46 : flight_46; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_129 = a_first & _a_first_T ? 7'h2f == auto_in_a_bits_source | flight_47 : flight_47; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_130 = a_first & _a_first_T ? 7'h30 == auto_in_a_bits_source | flight_48 : flight_48; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_131 = a_first & _a_first_T ? 7'h31 == auto_in_a_bits_source | flight_49 : flight_49; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_132 = a_first & _a_first_T ? 7'h32 == auto_in_a_bits_source | flight_50 : flight_50; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_133 = a_first & _a_first_T ? 7'h33 == auto_in_a_bits_source | flight_51 : flight_51; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_134 = a_first & _a_first_T ? 7'h34 == auto_in_a_bits_source | flight_52 : flight_52; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_135 = a_first & _a_first_T ? 7'h35 == auto_in_a_bits_source | flight_53 : flight_53; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_136 = a_first & _a_first_T ? 7'h36 == auto_in_a_bits_source | flight_54 : flight_54; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_137 = a_first & _a_first_T ? 7'h37 == auto_in_a_bits_source | flight_55 : flight_55; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_138 = a_first & _a_first_T ? 7'h38 == auto_in_a_bits_source | flight_56 : flight_56; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_139 = a_first & _a_first_T ? 7'h39 == auto_in_a_bits_source | flight_57 : flight_57; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_140 = a_first & _a_first_T ? 7'h3a == auto_in_a_bits_source | flight_58 : flight_58; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_141 = a_first & _a_first_T ? 7'h3b == auto_in_a_bits_source | flight_59 : flight_59; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_142 = a_first & _a_first_T ? 7'h3c == auto_in_a_bits_source | flight_60 : flight_60; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_143 = a_first & _a_first_T ? 7'h3d == auto_in_a_bits_source | flight_61 : flight_61; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_144 = a_first & _a_first_T ? 7'h3e == auto_in_a_bits_source | flight_62 : flight_62; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_145 = a_first & _a_first_T ? 7'h3f == auto_in_a_bits_source | flight_63 : flight_63; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_146 = a_first & _a_first_T ? 7'h40 == auto_in_a_bits_source | flight_64 : flight_64; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_147 = a_first & _a_first_T ? 7'h41 == auto_in_a_bits_source | flight_65 : flight_65; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_148 = a_first & _a_first_T ? 7'h42 == auto_in_a_bits_source | flight_66 : flight_66; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_149 = a_first & _a_first_T ? 7'h43 == auto_in_a_bits_source | flight_67 : flight_67; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_150 = a_first & _a_first_T ? 7'h44 == auto_in_a_bits_source | flight_68 : flight_68; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_151 = a_first & _a_first_T ? 7'h45 == auto_in_a_bits_source | flight_69 : flight_69; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_152 = a_first & _a_first_T ? 7'h46 == auto_in_a_bits_source | flight_70 : flight_70; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_153 = a_first & _a_first_T ? 7'h47 == auto_in_a_bits_source | flight_71 : flight_71; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_154 = a_first & _a_first_T ? 7'h48 == auto_in_a_bits_source | flight_72 : flight_72; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_155 = a_first & _a_first_T ? 7'h49 == auto_in_a_bits_source | flight_73 : flight_73; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_156 = a_first & _a_first_T ? 7'h4a == auto_in_a_bits_source | flight_74 : flight_74; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_157 = a_first & _a_first_T ? 7'h4b == auto_in_a_bits_source | flight_75 : flight_75; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_158 = a_first & _a_first_T ? 7'h4c == auto_in_a_bits_source | flight_76 : flight_76; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_159 = a_first & _a_first_T ? 7'h4d == auto_in_a_bits_source | flight_77 : flight_77; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_160 = a_first & _a_first_T ? 7'h4e == auto_in_a_bits_source | flight_78 : flight_78; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_161 = a_first & _a_first_T ? 7'h4f == auto_in_a_bits_source | flight_79 : flight_79; // @[FIFOFixer.scala 71:27 72:37]
  wire  _stalls_id_T_1 = _a_first_T & stalls_a_sel; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_5 = _a_first_T & stalls_a_sel_1; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_9 = _a_first_T & stalls_a_sel_2; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_13 = _a_first_T & stalls_a_sel_3; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_17 = _a_first_T & stalls_a_sel_4; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_21 = _a_first_T & stalls_a_sel_5; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_25 = _a_first_T & stalls_a_sel_6; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_29 = _a_first_T & stalls_a_sel_7; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_33 = _a_first_T & stalls_a_sel_8; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_37 = _a_first_T & stalls_a_sel_9; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_41 = _a_first_T & stalls_a_sel_10; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_45 = _a_first_T & stalls_a_sel_11; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_49 = _a_first_T & stalls_a_sel_12; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_53 = _a_first_T & stalls_a_sel_13; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_57 = _a_first_T & stalls_a_sel_14; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_61 = _a_first_T & stalls_a_sel_15; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_65 = _a_first_T & stalls_a_sel_16; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_69 = _a_first_T & stalls_a_sel_17; // @[FIFOFixer.scala 77:49]
  reg [19:0] TLFIFOFixer_3_covState; // @[Register tracking TLFIFOFixer_3 state]
  reg  TLFIFOFixer_3_covMap [0:1048575]; // @[Coverage map for TLFIFOFixer_3]
  wire  TLFIFOFixer_3_covMap_read_en; // @[Coverage map for TLFIFOFixer_3]
  wire [19:0] TLFIFOFixer_3_covMap_read_addr; // @[Coverage map for TLFIFOFixer_3]
  wire  TLFIFOFixer_3_covMap_read_data; // @[Coverage map for TLFIFOFixer_3]
  wire  TLFIFOFixer_3_covMap_write_data; // @[Coverage map for TLFIFOFixer_3]
  wire [19:0] TLFIFOFixer_3_covMap_write_addr; // @[Coverage map for TLFIFOFixer_3]
  wire  TLFIFOFixer_3_covMap_write_mask; // @[Coverage map for TLFIFOFixer_3]
  wire  TLFIFOFixer_3_covMap_write_en; // @[Coverage map for TLFIFOFixer_3]
  reg [29:0] TLFIFOFixer_3_covSum; // @[Sum of coverage map]
  wire [10:0] stalls_id_10_shl;
  wire [19:0] stalls_id_10_pad;
  wire [6:0] flight_77_shl;
  wire [19:0] flight_77_pad;
  wire [3:0] stalls_id_14_shl;
  wire [19:0] stalls_id_14_pad;
  wire [11:0] flight_41_shl;
  wire [19:0] flight_41_pad;
  wire [10:0] flight_53_shl;
  wire [19:0] flight_53_pad;
  wire [2:0] stalls_id_15_shl;
  wire [19:0] stalls_id_15_pad;
  wire [14:0] flight_1_shl;
  wire [19:0] flight_1_pad;
  wire [3:0] flight_40_shl;
  wire [19:0] flight_40_pad;
  wire [7:0] flight_23_shl;
  wire [19:0] flight_23_pad;
  wire [8:0] flight_72_shl;
  wire [19:0] flight_72_pad;
  wire [2:0] flight_34_shl;
  wire [19:0] flight_34_pad;
  wire [2:0] flight_47_shl;
  wire [19:0] flight_47_pad;
  wire [9:0] flight_56_shl;
  wire [19:0] flight_56_pad;
  wire [9:0] stalls_id_5_shl;
  wire [19:0] stalls_id_5_pad;
  wire [17:0] flight_20_shl;
  wire [19:0] flight_20_pad;
  wire [4:0] flight_60_shl;
  wire [19:0] flight_60_pad;
  wire [17:0] flight_71_shl;
  wire [19:0] flight_71_pad;
  wire [3:0] stalls_id_6_shl;
  wire [19:0] stalls_id_6_pad;
  wire [3:0] flight_49_shl;
  wire [19:0] flight_49_pad;
  wire [16:0] stalls_id_4_shl;
  wire [19:0] stalls_id_4_pad;
  wire [19:0] flight_12_shl;
  wire [19:0] flight_12_pad;
  wire [7:0] flight_8_shl;
  wire [19:0] flight_8_pad;
  wire [13:0] stalls_id_shl;
  wire [19:0] stalls_id_pad;
  wire [14:0] flight_9_shl;
  wire [19:0] flight_9_pad;
  wire [18:0] flight_57_shl;
  wire [19:0] flight_57_pad;
  wire [1:0] flight_75_shl;
  wire [19:0] flight_75_pad;
  wire [3:0] flight_48_shl;
  wire [19:0] flight_48_pad;
  wire [7:0] flight_10_shl;
  wire [19:0] flight_10_pad;
  wire [1:0] flight_32_shl;
  wire [19:0] flight_32_pad;
  wire [19:0] flight_61_shl;
  wire [19:0] flight_61_pad;
  wire [12:0] flight_5_shl;
  wire [19:0] flight_5_pad;
  wire  flight_39_shl;
  wire [19:0] flight_39_pad;
  wire [1:0] flight_19_shl;
  wire [19:0] flight_19_pad;
  wire [18:0] flight_58_shl;
  wire [19:0] flight_58_pad;
  wire [17:0] stalls_id_7_shl;
  wire [19:0] stalls_id_7_pad;
  wire [19:0] flight_73_shl;
  wire [19:0] flight_73_pad;
  wire [8:0] flight_21_shl;
  wire [19:0] flight_21_pad;
  wire [14:0] flight_62_shl;
  wire [19:0] flight_62_pad;
  wire [14:0] flight_76_shl;
  wire [19:0] flight_76_pad;
  wire [17:0] flight_15_shl;
  wire [19:0] flight_15_pad;
  wire [16:0] flight_14_shl;
  wire [19:0] flight_14_pad;
  wire [18:0] flight_51_shl;
  wire [19:0] flight_51_pad;
  wire [7:0] flight_37_shl;
  wire [19:0] flight_37_pad;
  wire [13:0] stalls_id_12_shl;
  wire [19:0] stalls_id_12_pad;
  wire [6:0] stalls_id_16_shl;
  wire [19:0] stalls_id_16_pad;
  wire [11:0] flight_13_shl;
  wire [19:0] flight_13_pad;
  wire [12:0] flight_78_shl;
  wire [19:0] flight_78_pad;
  wire [10:0] flight_46_shl;
  wire [19:0] flight_46_pad;
  wire [11:0] flight_74_shl;
  wire [19:0] flight_74_pad;
  wire [5:0] flight_16_shl;
  wire [19:0] flight_16_pad;
  wire [16:0] stalls_id_3_shl;
  wire [19:0] stalls_id_3_pad;
  wire [3:0] stalls_id_9_shl;
  wire [19:0] stalls_id_9_pad;
  wire [5:0] flight_7_shl;
  wire [19:0] flight_7_pad;
  wire [10:0] flight_69_shl;
  wire [19:0] flight_69_pad;
  wire [2:0] flight_79_shl;
  wire [19:0] flight_79_pad;
  wire [18:0] flight_0_shl;
  wire [19:0] flight_0_pad;
  wire [12:0] flight_38_shl;
  wire [19:0] flight_38_pad;
  wire  flight_30_shl;
  wire [19:0] flight_30_pad;
  wire [13:0] flight_22_shl;
  wire [19:0] flight_22_pad;
  wire [14:0] flight_59_shl;
  wire [19:0] flight_59_pad;
  wire [6:0] stalls_id_11_shl;
  wire [19:0] stalls_id_11_pad;
  wire [10:0] flight_55_shl;
  wire [19:0] flight_55_pad;
  wire [11:0] flight_67_shl;
  wire [19:0] flight_67_pad;
  wire [6:0] stalls_id_8_shl;
  wire [19:0] stalls_id_8_pad;
  wire [6:0] flight_65_shl;
  wire [19:0] flight_65_pad;
  wire [11:0] stalls_id_2_shl;
  wire [19:0] stalls_id_2_pad;
  wire [17:0] flight_64_shl;
  wire [19:0] flight_64_pad;
  wire [10:0] flight_45_shl;
  wire [19:0] flight_45_pad;
  wire [5:0] flight_11_shl;
  wire [19:0] flight_11_pad;
  wire [10:0] flight_6_shl;
  wire [19:0] flight_6_pad;
  wire [19:0] stalls_id_1_shl;
  wire [19:0] stalls_id_1_pad;
  wire [13:0] stalls_id_13_shl;
  wire [19:0] stalls_id_13_pad;
  wire [1:0] flight_31_shl;
  wire [19:0] flight_31_pad;
  wire [6:0] flight_66_shl;
  wire [19:0] flight_66_pad;
  wire [7:0] flight_70_shl;
  wire [19:0] flight_70_pad;
  wire [12:0] flight_3_shl;
  wire [19:0] flight_3_pad;
  wire [8:0] flight_42_shl;
  wire [19:0] flight_42_pad;
  wire [6:0] flight_25_shl;
  wire [19:0] flight_25_pad;
  wire  flight_17_shl;
  wire [19:0] flight_17_pad;
  wire [10:0] flight_36_shl;
  wire [19:0] flight_36_pad;
  wire [11:0] flight_2_shl;
  wire [19:0] flight_2_pad;
  wire [10:0] flight_29_shl;
  wire [19:0] flight_29_pad;
  wire [6:0] flight_27_shl;
  wire [19:0] flight_27_pad;
  wire  flight_33_shl;
  wire [19:0] flight_33_pad;
  wire [10:0] flight_35_shl;
  wire [19:0] flight_35_pad;
  wire [6:0] flight_68_shl;
  wire [19:0] flight_68_pad;
  wire [14:0] flight_4_shl;
  wire [19:0] flight_4_pad;
  wire [14:0] flight_28_shl;
  wire [19:0] flight_28_pad;
  wire [13:0] flight_18_shl;
  wire [19:0] flight_18_pad;
  wire [6:0] flight_63_shl;
  wire [19:0] flight_63_pad;
  wire [8:0] stalls_id_17_shl;
  wire [19:0] stalls_id_17_pad;
  wire [19:0] flight_54_shl;
  wire [19:0] flight_54_pad;
  wire [2:0] flight_50_shl;
  wire [19:0] flight_50_pad;
  wire [19:0] flight_44_shl;
  wire [19:0] flight_44_pad;
  wire [4:0] flight_43_shl;
  wire [19:0] flight_43_pad;
  wire [17:0] flight_52_shl;
  wire [19:0] flight_52_pad;
  wire [18:0] flight_26_shl;
  wire [19:0] flight_26_pad;
  wire  flight_24_shl;
  wire [19:0] flight_24_pad;
  wire [19:0] TLFIFOFixer_3_xor64;
  wire [19:0] TLFIFOFixer_3_xor31;
  wire [19:0] TLFIFOFixer_3_xor66;
  wire [19:0] TLFIFOFixer_3_xor32;
  wire [19:0] TLFIFOFixer_3_xor15;
  wire [19:0] TLFIFOFixer_3_xor68;
  wire [19:0] TLFIFOFixer_3_xor33;
  wire [19:0] TLFIFOFixer_3_xor70;
  wire [19:0] TLFIFOFixer_3_xor34;
  wire [19:0] TLFIFOFixer_3_xor16;
  wire [19:0] TLFIFOFixer_3_xor7;
  wire [19:0] TLFIFOFixer_3_xor72;
  wire [19:0] TLFIFOFixer_3_xor35;
  wire [19:0] TLFIFOFixer_3_xor74;
  wire [19:0] TLFIFOFixer_3_xor36;
  wire [19:0] TLFIFOFixer_3_xor17;
  wire [19:0] TLFIFOFixer_3_xor76;
  wire [19:0] TLFIFOFixer_3_xor37;
  wire [19:0] TLFIFOFixer_3_xor78;
  wire [19:0] TLFIFOFixer_3_xor38;
  wire [19:0] TLFIFOFixer_3_xor18;
  wire [19:0] TLFIFOFixer_3_xor8;
  wire [19:0] TLFIFOFixer_3_xor3;
  wire [19:0] TLFIFOFixer_3_xor80;
  wire [19:0] TLFIFOFixer_3_xor39;
  wire [19:0] TLFIFOFixer_3_xor82;
  wire [19:0] TLFIFOFixer_3_xor40;
  wire [19:0] TLFIFOFixer_3_xor19;
  wire [19:0] TLFIFOFixer_3_xor84;
  wire [19:0] TLFIFOFixer_3_xor41;
  wire [19:0] TLFIFOFixer_3_xor86;
  wire [19:0] TLFIFOFixer_3_xor42;
  wire [19:0] TLFIFOFixer_3_xor20;
  wire [19:0] TLFIFOFixer_3_xor9;
  wire [19:0] TLFIFOFixer_3_xor88;
  wire [19:0] TLFIFOFixer_3_xor43;
  wire [19:0] TLFIFOFixer_3_xor90;
  wire [19:0] TLFIFOFixer_3_xor44;
  wire [19:0] TLFIFOFixer_3_xor21;
  wire [19:0] TLFIFOFixer_3_xor92;
  wire [19:0] TLFIFOFixer_3_xor45;
  wire [19:0] TLFIFOFixer_3_xor93;
  wire [19:0] TLFIFOFixer_3_xor94;
  wire [19:0] TLFIFOFixer_3_xor46;
  wire [19:0] TLFIFOFixer_3_xor22;
  wire [19:0] TLFIFOFixer_3_xor10;
  wire [19:0] TLFIFOFixer_3_xor4;
  wire [19:0] TLFIFOFixer_3_xor1;
  wire [19:0] TLFIFOFixer_3_xor96;
  wire [19:0] TLFIFOFixer_3_xor47;
  wire [19:0] TLFIFOFixer_3_xor98;
  wire [19:0] TLFIFOFixer_3_xor48;
  wire [19:0] TLFIFOFixer_3_xor23;
  wire [19:0] TLFIFOFixer_3_xor100;
  wire [19:0] TLFIFOFixer_3_xor49;
  wire [19:0] TLFIFOFixer_3_xor102;
  wire [19:0] TLFIFOFixer_3_xor50;
  wire [19:0] TLFIFOFixer_3_xor24;
  wire [19:0] TLFIFOFixer_3_xor11;
  wire [19:0] TLFIFOFixer_3_xor104;
  wire [19:0] TLFIFOFixer_3_xor51;
  wire [19:0] TLFIFOFixer_3_xor106;
  wire [19:0] TLFIFOFixer_3_xor52;
  wire [19:0] TLFIFOFixer_3_xor25;
  wire [19:0] TLFIFOFixer_3_xor108;
  wire [19:0] TLFIFOFixer_3_xor53;
  wire [19:0] TLFIFOFixer_3_xor110;
  wire [19:0] TLFIFOFixer_3_xor54;
  wire [19:0] TLFIFOFixer_3_xor26;
  wire [19:0] TLFIFOFixer_3_xor12;
  wire [19:0] TLFIFOFixer_3_xor5;
  wire [19:0] TLFIFOFixer_3_xor112;
  wire [19:0] TLFIFOFixer_3_xor55;
  wire [19:0] TLFIFOFixer_3_xor114;
  wire [19:0] TLFIFOFixer_3_xor56;
  wire [19:0] TLFIFOFixer_3_xor27;
  wire [19:0] TLFIFOFixer_3_xor116;
  wire [19:0] TLFIFOFixer_3_xor57;
  wire [19:0] TLFIFOFixer_3_xor118;
  wire [19:0] TLFIFOFixer_3_xor58;
  wire [19:0] TLFIFOFixer_3_xor28;
  wire [19:0] TLFIFOFixer_3_xor13;
  wire [19:0] TLFIFOFixer_3_xor120;
  wire [19:0] TLFIFOFixer_3_xor59;
  wire [19:0] TLFIFOFixer_3_xor122;
  wire [19:0] TLFIFOFixer_3_xor60;
  wire [19:0] TLFIFOFixer_3_xor29;
  wire [19:0] TLFIFOFixer_3_xor124;
  wire [19:0] TLFIFOFixer_3_xor61;
  wire [19:0] TLFIFOFixer_3_xor125;
  wire [19:0] TLFIFOFixer_3_xor126;
  wire [19:0] TLFIFOFixer_3_xor62;
  wire [19:0] TLFIFOFixer_3_xor30;
  wire [19:0] TLFIFOFixer_3_xor14;
  wire [19:0] TLFIFOFixer_3_xor6;
  wire [19:0] TLFIFOFixer_3_xor2;
  wire [19:0] TLFIFOFixer_3_xor0;
  assign auto_in_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  assign auto_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = auto_in_a_valid & _bundleIn_0_a_ready_T; // @[FIFOFixer.scala 87:33]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLFIFOFixer_3_covMap_read_en = 1'h1;
  assign TLFIFOFixer_3_covMap_read_addr = TLFIFOFixer_3_covState;
  assign TLFIFOFixer_3_covMap_read_data = TLFIFOFixer_3_covMap[TLFIFOFixer_3_covMap_read_addr]; // @[Coverage map for TLFIFOFixer_3]
  assign TLFIFOFixer_3_covMap_write_data = 1'h1;
  assign TLFIFOFixer_3_covMap_write_addr = TLFIFOFixer_3_covState;
  assign TLFIFOFixer_3_covMap_write_mask = 1'h1;
  assign TLFIFOFixer_3_covMap_write_en = ~metaReset;
  assign stalls_id_10_shl = {stalls_id_10, 8'h0};
  assign stalls_id_10_pad = {9'h0,stalls_id_10_shl};
  assign flight_77_shl = {flight_77, 6'h0};
  assign flight_77_pad = {13'h0,flight_77_shl};
  assign stalls_id_14_shl = {stalls_id_14, 1'h0};
  assign stalls_id_14_pad = {16'h0,stalls_id_14_shl};
  assign flight_41_shl = {flight_41, 11'h0};
  assign flight_41_pad = {8'h0,flight_41_shl};
  assign flight_53_shl = {flight_53, 10'h0};
  assign flight_53_pad = {9'h0,flight_53_shl};
  assign stalls_id_15_shl = stalls_id_15;
  assign stalls_id_15_pad = {17'h0,stalls_id_15_shl};
  assign flight_1_shl = {flight_1, 14'h0};
  assign flight_1_pad = {5'h0,flight_1_shl};
  assign flight_40_shl = {flight_40, 3'h0};
  assign flight_40_pad = {16'h0,flight_40_shl};
  assign flight_23_shl = {flight_23, 7'h0};
  assign flight_23_pad = {12'h0,flight_23_shl};
  assign flight_72_shl = {flight_72, 8'h0};
  assign flight_72_pad = {11'h0,flight_72_shl};
  assign flight_34_shl = {flight_34, 2'h0};
  assign flight_34_pad = {17'h0,flight_34_shl};
  assign flight_47_shl = {flight_47, 2'h0};
  assign flight_47_pad = {17'h0,flight_47_shl};
  assign flight_56_shl = {flight_56, 9'h0};
  assign flight_56_pad = {10'h0,flight_56_shl};
  assign stalls_id_5_shl = {stalls_id_5, 7'h0};
  assign stalls_id_5_pad = {10'h0,stalls_id_5_shl};
  assign flight_20_shl = {flight_20, 17'h0};
  assign flight_20_pad = {2'h0,flight_20_shl};
  assign flight_60_shl = {flight_60, 4'h0};
  assign flight_60_pad = {15'h0,flight_60_shl};
  assign flight_71_shl = {flight_71, 17'h0};
  assign flight_71_pad = {2'h0,flight_71_shl};
  assign stalls_id_6_shl = {stalls_id_6, 1'h0};
  assign stalls_id_6_pad = {16'h0,stalls_id_6_shl};
  assign flight_49_shl = {flight_49, 3'h0};
  assign flight_49_pad = {16'h0,flight_49_shl};
  assign stalls_id_4_shl = {stalls_id_4, 14'h0};
  assign stalls_id_4_pad = {3'h0,stalls_id_4_shl};
  assign flight_12_shl = {flight_12, 19'h0};
  assign flight_12_pad = flight_12_shl;
  assign flight_8_shl = {flight_8, 7'h0};
  assign flight_8_pad = {12'h0,flight_8_shl};
  assign stalls_id_shl = {stalls_id, 11'h0};
  assign stalls_id_pad = {6'h0,stalls_id_shl};
  assign flight_9_shl = {flight_9, 14'h0};
  assign flight_9_pad = {5'h0,flight_9_shl};
  assign flight_57_shl = {flight_57, 18'h0};
  assign flight_57_pad = {1'h0,flight_57_shl};
  assign flight_75_shl = {flight_75, 1'h0};
  assign flight_75_pad = {18'h0,flight_75_shl};
  assign flight_48_shl = {flight_48, 3'h0};
  assign flight_48_pad = {16'h0,flight_48_shl};
  assign flight_10_shl = {flight_10, 7'h0};
  assign flight_10_pad = {12'h0,flight_10_shl};
  assign flight_32_shl = {flight_32, 1'h0};
  assign flight_32_pad = {18'h0,flight_32_shl};
  assign flight_61_shl = {flight_61, 19'h0};
  assign flight_61_pad = flight_61_shl;
  assign flight_5_shl = {flight_5, 12'h0};
  assign flight_5_pad = {7'h0,flight_5_shl};
  assign flight_39_shl = flight_39;
  assign flight_39_pad = {19'h0,flight_39_shl};
  assign flight_19_shl = {flight_19, 1'h0};
  assign flight_19_pad = {18'h0,flight_19_shl};
  assign flight_58_shl = {flight_58, 18'h0};
  assign flight_58_pad = {1'h0,flight_58_shl};
  assign stalls_id_7_shl = {stalls_id_7, 15'h0};
  assign stalls_id_7_pad = {2'h0,stalls_id_7_shl};
  assign flight_73_shl = {flight_73, 19'h0};
  assign flight_73_pad = flight_73_shl;
  assign flight_21_shl = {flight_21, 8'h0};
  assign flight_21_pad = {11'h0,flight_21_shl};
  assign flight_62_shl = {flight_62, 14'h0};
  assign flight_62_pad = {5'h0,flight_62_shl};
  assign flight_76_shl = {flight_76, 14'h0};
  assign flight_76_pad = {5'h0,flight_76_shl};
  assign flight_15_shl = {flight_15, 17'h0};
  assign flight_15_pad = {2'h0,flight_15_shl};
  assign flight_14_shl = {flight_14, 16'h0};
  assign flight_14_pad = {3'h0,flight_14_shl};
  assign flight_51_shl = {flight_51, 18'h0};
  assign flight_51_pad = {1'h0,flight_51_shl};
  assign flight_37_shl = {flight_37, 7'h0};
  assign flight_37_pad = {12'h0,flight_37_shl};
  assign stalls_id_12_shl = {stalls_id_12, 11'h0};
  assign stalls_id_12_pad = {6'h0,stalls_id_12_shl};
  assign stalls_id_16_shl = {stalls_id_16, 4'h0};
  assign stalls_id_16_pad = {13'h0,stalls_id_16_shl};
  assign flight_13_shl = {flight_13, 11'h0};
  assign flight_13_pad = {8'h0,flight_13_shl};
  assign flight_78_shl = {flight_78, 12'h0};
  assign flight_78_pad = {7'h0,flight_78_shl};
  assign flight_46_shl = {flight_46, 10'h0};
  assign flight_46_pad = {9'h0,flight_46_shl};
  assign flight_74_shl = {flight_74, 11'h0};
  assign flight_74_pad = {8'h0,flight_74_shl};
  assign flight_16_shl = {flight_16, 5'h0};
  assign flight_16_pad = {14'h0,flight_16_shl};
  assign stalls_id_3_shl = {stalls_id_3, 14'h0};
  assign stalls_id_3_pad = {3'h0,stalls_id_3_shl};
  assign stalls_id_9_shl = {stalls_id_9, 1'h0};
  assign stalls_id_9_pad = {16'h0,stalls_id_9_shl};
  assign flight_7_shl = {flight_7, 5'h0};
  assign flight_7_pad = {14'h0,flight_7_shl};
  assign flight_69_shl = {flight_69, 10'h0};
  assign flight_69_pad = {9'h0,flight_69_shl};
  assign flight_79_shl = {flight_79, 2'h0};
  assign flight_79_pad = {17'h0,flight_79_shl};
  assign flight_0_shl = {flight_0, 18'h0};
  assign flight_0_pad = {1'h0,flight_0_shl};
  assign flight_38_shl = {flight_38, 12'h0};
  assign flight_38_pad = {7'h0,flight_38_shl};
  assign flight_30_shl = flight_30;
  assign flight_30_pad = {19'h0,flight_30_shl};
  assign flight_22_shl = {flight_22, 13'h0};
  assign flight_22_pad = {6'h0,flight_22_shl};
  assign flight_59_shl = {flight_59, 14'h0};
  assign flight_59_pad = {5'h0,flight_59_shl};
  assign stalls_id_11_shl = {stalls_id_11, 4'h0};
  assign stalls_id_11_pad = {13'h0,stalls_id_11_shl};
  assign flight_55_shl = {flight_55, 10'h0};
  assign flight_55_pad = {9'h0,flight_55_shl};
  assign flight_67_shl = {flight_67, 11'h0};
  assign flight_67_pad = {8'h0,flight_67_shl};
  assign stalls_id_8_shl = {stalls_id_8, 4'h0};
  assign stalls_id_8_pad = {13'h0,stalls_id_8_shl};
  assign flight_65_shl = {flight_65, 6'h0};
  assign flight_65_pad = {13'h0,flight_65_shl};
  assign stalls_id_2_shl = {stalls_id_2, 9'h0};
  assign stalls_id_2_pad = {8'h0,stalls_id_2_shl};
  assign flight_64_shl = {flight_64, 17'h0};
  assign flight_64_pad = {2'h0,flight_64_shl};
  assign flight_45_shl = {flight_45, 10'h0};
  assign flight_45_pad = {9'h0,flight_45_shl};
  assign flight_11_shl = {flight_11, 5'h0};
  assign flight_11_pad = {14'h0,flight_11_shl};
  assign flight_6_shl = {flight_6, 10'h0};
  assign flight_6_pad = {9'h0,flight_6_shl};
  assign stalls_id_1_shl = {stalls_id_1, 17'h0};
  assign stalls_id_1_pad = stalls_id_1_shl;
  assign stalls_id_13_shl = {stalls_id_13, 11'h0};
  assign stalls_id_13_pad = {6'h0,stalls_id_13_shl};
  assign flight_31_shl = {flight_31, 1'h0};
  assign flight_31_pad = {18'h0,flight_31_shl};
  assign flight_66_shl = {flight_66, 6'h0};
  assign flight_66_pad = {13'h0,flight_66_shl};
  assign flight_70_shl = {flight_70, 7'h0};
  assign flight_70_pad = {12'h0,flight_70_shl};
  assign flight_3_shl = {flight_3, 12'h0};
  assign flight_3_pad = {7'h0,flight_3_shl};
  assign flight_42_shl = {flight_42, 8'h0};
  assign flight_42_pad = {11'h0,flight_42_shl};
  assign flight_25_shl = {flight_25, 6'h0};
  assign flight_25_pad = {13'h0,flight_25_shl};
  assign flight_17_shl = flight_17;
  assign flight_17_pad = {19'h0,flight_17_shl};
  assign flight_36_shl = {flight_36, 10'h0};
  assign flight_36_pad = {9'h0,flight_36_shl};
  assign flight_2_shl = {flight_2, 11'h0};
  assign flight_2_pad = {8'h0,flight_2_shl};
  assign flight_29_shl = {flight_29, 10'h0};
  assign flight_29_pad = {9'h0,flight_29_shl};
  assign flight_27_shl = {flight_27, 6'h0};
  assign flight_27_pad = {13'h0,flight_27_shl};
  assign flight_33_shl = flight_33;
  assign flight_33_pad = {19'h0,flight_33_shl};
  assign flight_35_shl = {flight_35, 10'h0};
  assign flight_35_pad = {9'h0,flight_35_shl};
  assign flight_68_shl = {flight_68, 6'h0};
  assign flight_68_pad = {13'h0,flight_68_shl};
  assign flight_4_shl = {flight_4, 14'h0};
  assign flight_4_pad = {5'h0,flight_4_shl};
  assign flight_28_shl = {flight_28, 14'h0};
  assign flight_28_pad = {5'h0,flight_28_shl};
  assign flight_18_shl = {flight_18, 13'h0};
  assign flight_18_pad = {6'h0,flight_18_shl};
  assign flight_63_shl = {flight_63, 6'h0};
  assign flight_63_pad = {13'h0,flight_63_shl};
  assign stalls_id_17_shl = {stalls_id_17, 6'h0};
  assign stalls_id_17_pad = {11'h0,stalls_id_17_shl};
  assign flight_54_shl = {flight_54, 19'h0};
  assign flight_54_pad = flight_54_shl;
  assign flight_50_shl = {flight_50, 2'h0};
  assign flight_50_pad = {17'h0,flight_50_shl};
  assign flight_44_shl = {flight_44, 19'h0};
  assign flight_44_pad = flight_44_shl;
  assign flight_43_shl = {flight_43, 4'h0};
  assign flight_43_pad = {15'h0,flight_43_shl};
  assign flight_52_shl = {flight_52, 17'h0};
  assign flight_52_pad = {2'h0,flight_52_shl};
  assign flight_26_shl = {flight_26, 18'h0};
  assign flight_26_pad = {1'h0,flight_26_shl};
  assign flight_24_shl = flight_24;
  assign flight_24_pad = {19'h0,flight_24_shl};
  assign TLFIFOFixer_3_xor64 = flight_77_pad ^ stalls_id_14_pad;
  assign TLFIFOFixer_3_xor31 = stalls_id_10_pad ^ TLFIFOFixer_3_xor64;
  assign TLFIFOFixer_3_xor66 = flight_53_pad ^ stalls_id_15_pad;
  assign TLFIFOFixer_3_xor32 = flight_41_pad ^ TLFIFOFixer_3_xor66;
  assign TLFIFOFixer_3_xor15 = TLFIFOFixer_3_xor31 ^ TLFIFOFixer_3_xor32;
  assign TLFIFOFixer_3_xor68 = flight_40_pad ^ flight_23_pad;
  assign TLFIFOFixer_3_xor33 = flight_1_pad ^ TLFIFOFixer_3_xor68;
  assign TLFIFOFixer_3_xor70 = flight_34_pad ^ flight_47_pad;
  assign TLFIFOFixer_3_xor34 = flight_72_pad ^ TLFIFOFixer_3_xor70;
  assign TLFIFOFixer_3_xor16 = TLFIFOFixer_3_xor33 ^ TLFIFOFixer_3_xor34;
  assign TLFIFOFixer_3_xor7 = TLFIFOFixer_3_xor15 ^ TLFIFOFixer_3_xor16;
  assign TLFIFOFixer_3_xor72 = stalls_id_5_pad ^ flight_20_pad;
  assign TLFIFOFixer_3_xor35 = flight_56_pad ^ TLFIFOFixer_3_xor72;
  assign TLFIFOFixer_3_xor74 = flight_71_pad ^ stalls_id_6_pad;
  assign TLFIFOFixer_3_xor36 = flight_60_pad ^ TLFIFOFixer_3_xor74;
  assign TLFIFOFixer_3_xor17 = TLFIFOFixer_3_xor35 ^ TLFIFOFixer_3_xor36;
  assign TLFIFOFixer_3_xor76 = stalls_id_4_pad ^ flight_12_pad;
  assign TLFIFOFixer_3_xor37 = flight_49_pad ^ TLFIFOFixer_3_xor76;
  assign TLFIFOFixer_3_xor78 = stalls_id_pad ^ flight_9_pad;
  assign TLFIFOFixer_3_xor38 = flight_8_pad ^ TLFIFOFixer_3_xor78;
  assign TLFIFOFixer_3_xor18 = TLFIFOFixer_3_xor37 ^ TLFIFOFixer_3_xor38;
  assign TLFIFOFixer_3_xor8 = TLFIFOFixer_3_xor17 ^ TLFIFOFixer_3_xor18;
  assign TLFIFOFixer_3_xor3 = TLFIFOFixer_3_xor7 ^ TLFIFOFixer_3_xor8;
  assign TLFIFOFixer_3_xor80 = flight_75_pad ^ flight_48_pad;
  assign TLFIFOFixer_3_xor39 = flight_57_pad ^ TLFIFOFixer_3_xor80;
  assign TLFIFOFixer_3_xor82 = flight_32_pad ^ flight_61_pad;
  assign TLFIFOFixer_3_xor40 = flight_10_pad ^ TLFIFOFixer_3_xor82;
  assign TLFIFOFixer_3_xor19 = TLFIFOFixer_3_xor39 ^ TLFIFOFixer_3_xor40;
  assign TLFIFOFixer_3_xor84 = flight_39_pad ^ flight_19_pad;
  assign TLFIFOFixer_3_xor41 = flight_5_pad ^ TLFIFOFixer_3_xor84;
  assign TLFIFOFixer_3_xor86 = stalls_id_7_pad ^ flight_73_pad;
  assign TLFIFOFixer_3_xor42 = flight_58_pad ^ TLFIFOFixer_3_xor86;
  assign TLFIFOFixer_3_xor20 = TLFIFOFixer_3_xor41 ^ TLFIFOFixer_3_xor42;
  assign TLFIFOFixer_3_xor9 = TLFIFOFixer_3_xor19 ^ TLFIFOFixer_3_xor20;
  assign TLFIFOFixer_3_xor88 = flight_62_pad ^ flight_76_pad;
  assign TLFIFOFixer_3_xor43 = flight_21_pad ^ TLFIFOFixer_3_xor88;
  assign TLFIFOFixer_3_xor90 = flight_14_pad ^ flight_51_pad;
  assign TLFIFOFixer_3_xor44 = flight_15_pad ^ TLFIFOFixer_3_xor90;
  assign TLFIFOFixer_3_xor21 = TLFIFOFixer_3_xor43 ^ TLFIFOFixer_3_xor44;
  assign TLFIFOFixer_3_xor92 = stalls_id_12_pad ^ stalls_id_16_pad;
  assign TLFIFOFixer_3_xor45 = flight_37_pad ^ TLFIFOFixer_3_xor92;
  assign TLFIFOFixer_3_xor93 = flight_13_pad ^ flight_78_pad;
  assign TLFIFOFixer_3_xor94 = flight_46_pad ^ flight_74_pad;
  assign TLFIFOFixer_3_xor46 = TLFIFOFixer_3_xor93 ^ TLFIFOFixer_3_xor94;
  assign TLFIFOFixer_3_xor22 = TLFIFOFixer_3_xor45 ^ TLFIFOFixer_3_xor46;
  assign TLFIFOFixer_3_xor10 = TLFIFOFixer_3_xor21 ^ TLFIFOFixer_3_xor22;
  assign TLFIFOFixer_3_xor4 = TLFIFOFixer_3_xor9 ^ TLFIFOFixer_3_xor10;
  assign TLFIFOFixer_3_xor1 = TLFIFOFixer_3_xor3 ^ TLFIFOFixer_3_xor4;
  assign TLFIFOFixer_3_xor96 = stalls_id_3_pad ^ stalls_id_9_pad;
  assign TLFIFOFixer_3_xor47 = flight_16_pad ^ TLFIFOFixer_3_xor96;
  assign TLFIFOFixer_3_xor98 = flight_69_pad ^ flight_79_pad;
  assign TLFIFOFixer_3_xor48 = flight_7_pad ^ TLFIFOFixer_3_xor98;
  assign TLFIFOFixer_3_xor23 = TLFIFOFixer_3_xor47 ^ TLFIFOFixer_3_xor48;
  assign TLFIFOFixer_3_xor100 = flight_38_pad ^ flight_30_pad;
  assign TLFIFOFixer_3_xor49 = flight_0_pad ^ TLFIFOFixer_3_xor100;
  assign TLFIFOFixer_3_xor102 = flight_59_pad ^ stalls_id_11_pad;
  assign TLFIFOFixer_3_xor50 = flight_22_pad ^ TLFIFOFixer_3_xor102;
  assign TLFIFOFixer_3_xor24 = TLFIFOFixer_3_xor49 ^ TLFIFOFixer_3_xor50;
  assign TLFIFOFixer_3_xor11 = TLFIFOFixer_3_xor23 ^ TLFIFOFixer_3_xor24;
  assign TLFIFOFixer_3_xor104 = flight_67_pad ^ stalls_id_8_pad;
  assign TLFIFOFixer_3_xor51 = flight_55_pad ^ TLFIFOFixer_3_xor104;
  assign TLFIFOFixer_3_xor106 = stalls_id_2_pad ^ flight_64_pad;
  assign TLFIFOFixer_3_xor52 = flight_65_pad ^ TLFIFOFixer_3_xor106;
  assign TLFIFOFixer_3_xor25 = TLFIFOFixer_3_xor51 ^ TLFIFOFixer_3_xor52;
  assign TLFIFOFixer_3_xor108 = flight_11_pad ^ flight_6_pad;
  assign TLFIFOFixer_3_xor53 = flight_45_pad ^ TLFIFOFixer_3_xor108;
  assign TLFIFOFixer_3_xor110 = stalls_id_13_pad ^ flight_31_pad;
  assign TLFIFOFixer_3_xor54 = stalls_id_1_pad ^ TLFIFOFixer_3_xor110;
  assign TLFIFOFixer_3_xor26 = TLFIFOFixer_3_xor53 ^ TLFIFOFixer_3_xor54;
  assign TLFIFOFixer_3_xor12 = TLFIFOFixer_3_xor25 ^ TLFIFOFixer_3_xor26;
  assign TLFIFOFixer_3_xor5 = TLFIFOFixer_3_xor11 ^ TLFIFOFixer_3_xor12;
  assign TLFIFOFixer_3_xor112 = flight_70_pad ^ flight_3_pad;
  assign TLFIFOFixer_3_xor55 = flight_66_pad ^ TLFIFOFixer_3_xor112;
  assign TLFIFOFixer_3_xor114 = flight_25_pad ^ flight_17_pad;
  assign TLFIFOFixer_3_xor56 = flight_42_pad ^ TLFIFOFixer_3_xor114;
  assign TLFIFOFixer_3_xor27 = TLFIFOFixer_3_xor55 ^ TLFIFOFixer_3_xor56;
  assign TLFIFOFixer_3_xor116 = flight_2_pad ^ flight_29_pad;
  assign TLFIFOFixer_3_xor57 = flight_36_pad ^ TLFIFOFixer_3_xor116;
  assign TLFIFOFixer_3_xor118 = flight_33_pad ^ flight_35_pad;
  assign TLFIFOFixer_3_xor58 = flight_27_pad ^ TLFIFOFixer_3_xor118;
  assign TLFIFOFixer_3_xor28 = TLFIFOFixer_3_xor57 ^ TLFIFOFixer_3_xor58;
  assign TLFIFOFixer_3_xor13 = TLFIFOFixer_3_xor27 ^ TLFIFOFixer_3_xor28;
  assign TLFIFOFixer_3_xor120 = flight_4_pad ^ flight_28_pad;
  assign TLFIFOFixer_3_xor59 = flight_68_pad ^ TLFIFOFixer_3_xor120;
  assign TLFIFOFixer_3_xor122 = flight_63_pad ^ stalls_id_17_pad;
  assign TLFIFOFixer_3_xor60 = flight_18_pad ^ TLFIFOFixer_3_xor122;
  assign TLFIFOFixer_3_xor29 = TLFIFOFixer_3_xor59 ^ TLFIFOFixer_3_xor60;
  assign TLFIFOFixer_3_xor124 = flight_50_pad ^ flight_44_pad;
  assign TLFIFOFixer_3_xor61 = flight_54_pad ^ TLFIFOFixer_3_xor124;
  assign TLFIFOFixer_3_xor125 = flight_43_pad ^ flight_52_pad;
  assign TLFIFOFixer_3_xor126 = flight_26_pad ^ flight_24_pad;
  assign TLFIFOFixer_3_xor62 = TLFIFOFixer_3_xor125 ^ TLFIFOFixer_3_xor126;
  assign TLFIFOFixer_3_xor30 = TLFIFOFixer_3_xor61 ^ TLFIFOFixer_3_xor62;
  assign TLFIFOFixer_3_xor14 = TLFIFOFixer_3_xor29 ^ TLFIFOFixer_3_xor30;
  assign TLFIFOFixer_3_xor6 = TLFIFOFixer_3_xor13 ^ TLFIFOFixer_3_xor14;
  assign TLFIFOFixer_3_xor2 = TLFIFOFixer_3_xor5 ^ TLFIFOFixer_3_xor6;
  assign TLFIFOFixer_3_xor0 = TLFIFOFixer_3_xor1 ^ TLFIFOFixer_3_xor2;
  assign io_covSum = TLFIFOFixer_3_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin
      if (a_first) begin
        if (a_first_beats1_opdata) begin
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_64 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h40 == auto_out_d_bits_source) begin
        flight_64 <= 1'h0;
      end else begin
        flight_64 <= _GEN_146;
      end
    end else begin
      flight_64 <= _GEN_146;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_65 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h41 == auto_out_d_bits_source) begin
        flight_65 <= 1'h0;
      end else begin
        flight_65 <= _GEN_147;
      end
    end else begin
      flight_65 <= _GEN_147;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_66 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h42 == auto_out_d_bits_source) begin
        flight_66 <= 1'h0;
      end else begin
        flight_66 <= _GEN_148;
      end
    end else begin
      flight_66 <= _GEN_148;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_67 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h43 == auto_out_d_bits_source) begin
        flight_67 <= 1'h0;
      end else begin
        flight_67 <= _GEN_149;
      end
    end else begin
      flight_67 <= _GEN_149;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_68 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h44 == auto_out_d_bits_source) begin
        flight_68 <= 1'h0;
      end else begin
        flight_68 <= _GEN_150;
      end
    end else begin
      flight_68 <= _GEN_150;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_69 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h45 == auto_out_d_bits_source) begin
        flight_69 <= 1'h0;
      end else begin
        flight_69 <= _GEN_151;
      end
    end else begin
      flight_69 <= _GEN_151;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_70 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h46 == auto_out_d_bits_source) begin
        flight_70 <= 1'h0;
      end else begin
        flight_70 <= _GEN_152;
      end
    end else begin
      flight_70 <= _GEN_152;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_71 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h47 == auto_out_d_bits_source) begin
        flight_71 <= 1'h0;
      end else begin
        flight_71 <= _GEN_153;
      end
    end else begin
      flight_71 <= _GEN_153;
    end
    if (_stalls_id_T_1) begin // @[Reg.scala 17:18]
      stalls_id <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_72 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h48 == auto_out_d_bits_source) begin
        flight_72 <= 1'h0;
      end else begin
        flight_72 <= _GEN_154;
      end
    end else begin
      flight_72 <= _GEN_154;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_73 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h49 == auto_out_d_bits_source) begin
        flight_73 <= 1'h0;
      end else begin
        flight_73 <= _GEN_155;
      end
    end else begin
      flight_73 <= _GEN_155;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_74 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h4a == auto_out_d_bits_source) begin
        flight_74 <= 1'h0;
      end else begin
        flight_74 <= _GEN_156;
      end
    end else begin
      flight_74 <= _GEN_156;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_75 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h4b == auto_out_d_bits_source) begin
        flight_75 <= 1'h0;
      end else begin
        flight_75 <= _GEN_157;
      end
    end else begin
      flight_75 <= _GEN_157;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_76 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h4c == auto_out_d_bits_source) begin
        flight_76 <= 1'h0;
      end else begin
        flight_76 <= _GEN_158;
      end
    end else begin
      flight_76 <= _GEN_158;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_77 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h4d == auto_out_d_bits_source) begin
        flight_77 <= 1'h0;
      end else begin
        flight_77 <= _GEN_159;
      end
    end else begin
      flight_77 <= _GEN_159;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_78 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h4e == auto_out_d_bits_source) begin
        flight_78 <= 1'h0;
      end else begin
        flight_78 <= _GEN_160;
      end
    end else begin
      flight_78 <= _GEN_160;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_79 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h4f == auto_out_d_bits_source) begin
        flight_79 <= 1'h0;
      end else begin
        flight_79 <= _GEN_161;
      end
    end else begin
      flight_79 <= _GEN_161;
    end
    if (_stalls_id_T_5) begin // @[Reg.scala 17:18]
      stalls_id_1 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_0 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h0 == auto_out_d_bits_source) begin
        flight_0 <= 1'h0;
      end else begin
        flight_0 <= _GEN_82;
      end
    end else begin
      flight_0 <= _GEN_82;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_1 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h1 == auto_out_d_bits_source) begin
        flight_1 <= 1'h0;
      end else begin
        flight_1 <= _GEN_83;
      end
    end else begin
      flight_1 <= _GEN_83;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_2 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h2 == auto_out_d_bits_source) begin
        flight_2 <= 1'h0;
      end else begin
        flight_2 <= _GEN_84;
      end
    end else begin
      flight_2 <= _GEN_84;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_3 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h3 == auto_out_d_bits_source) begin
        flight_3 <= 1'h0;
      end else begin
        flight_3 <= _GEN_85;
      end
    end else begin
      flight_3 <= _GEN_85;
    end
    if (_stalls_id_T_9) begin // @[Reg.scala 17:18]
      stalls_id_2 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_4 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h4 == auto_out_d_bits_source) begin
        flight_4 <= 1'h0;
      end else begin
        flight_4 <= _GEN_86;
      end
    end else begin
      flight_4 <= _GEN_86;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_5 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h5 == auto_out_d_bits_source) begin
        flight_5 <= 1'h0;
      end else begin
        flight_5 <= _GEN_87;
      end
    end else begin
      flight_5 <= _GEN_87;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_6 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h6 == auto_out_d_bits_source) begin
        flight_6 <= 1'h0;
      end else begin
        flight_6 <= _GEN_88;
      end
    end else begin
      flight_6 <= _GEN_88;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_7 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h7 == auto_out_d_bits_source) begin
        flight_7 <= 1'h0;
      end else begin
        flight_7 <= _GEN_89;
      end
    end else begin
      flight_7 <= _GEN_89;
    end
    if (_stalls_id_T_13) begin // @[Reg.scala 17:18]
      stalls_id_3 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_8 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h8 == auto_out_d_bits_source) begin
        flight_8 <= 1'h0;
      end else begin
        flight_8 <= _GEN_90;
      end
    end else begin
      flight_8 <= _GEN_90;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_9 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h9 == auto_out_d_bits_source) begin
        flight_9 <= 1'h0;
      end else begin
        flight_9 <= _GEN_91;
      end
    end else begin
      flight_9 <= _GEN_91;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_10 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'ha == auto_out_d_bits_source) begin
        flight_10 <= 1'h0;
      end else begin
        flight_10 <= _GEN_92;
      end
    end else begin
      flight_10 <= _GEN_92;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_11 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'hb == auto_out_d_bits_source) begin
        flight_11 <= 1'h0;
      end else begin
        flight_11 <= _GEN_93;
      end
    end else begin
      flight_11 <= _GEN_93;
    end
    if (_stalls_id_T_17) begin // @[Reg.scala 17:18]
      stalls_id_4 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_12 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'hc == auto_out_d_bits_source) begin
        flight_12 <= 1'h0;
      end else begin
        flight_12 <= _GEN_94;
      end
    end else begin
      flight_12 <= _GEN_94;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_13 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'hd == auto_out_d_bits_source) begin
        flight_13 <= 1'h0;
      end else begin
        flight_13 <= _GEN_95;
      end
    end else begin
      flight_13 <= _GEN_95;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_14 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'he == auto_out_d_bits_source) begin
        flight_14 <= 1'h0;
      end else begin
        flight_14 <= _GEN_96;
      end
    end else begin
      flight_14 <= _GEN_96;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_15 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'hf == auto_out_d_bits_source) begin
        flight_15 <= 1'h0;
      end else begin
        flight_15 <= _GEN_97;
      end
    end else begin
      flight_15 <= _GEN_97;
    end
    if (_stalls_id_T_21) begin // @[Reg.scala 17:18]
      stalls_id_5 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_16 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h10 == auto_out_d_bits_source) begin
        flight_16 <= 1'h0;
      end else begin
        flight_16 <= _GEN_98;
      end
    end else begin
      flight_16 <= _GEN_98;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_17 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h11 == auto_out_d_bits_source) begin
        flight_17 <= 1'h0;
      end else begin
        flight_17 <= _GEN_99;
      end
    end else begin
      flight_17 <= _GEN_99;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_18 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h12 == auto_out_d_bits_source) begin
        flight_18 <= 1'h0;
      end else begin
        flight_18 <= _GEN_100;
      end
    end else begin
      flight_18 <= _GEN_100;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_19 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h13 == auto_out_d_bits_source) begin
        flight_19 <= 1'h0;
      end else begin
        flight_19 <= _GEN_101;
      end
    end else begin
      flight_19 <= _GEN_101;
    end
    if (_stalls_id_T_25) begin // @[Reg.scala 17:18]
      stalls_id_6 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_20 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h14 == auto_out_d_bits_source) begin
        flight_20 <= 1'h0;
      end else begin
        flight_20 <= _GEN_102;
      end
    end else begin
      flight_20 <= _GEN_102;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_21 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h15 == auto_out_d_bits_source) begin
        flight_21 <= 1'h0;
      end else begin
        flight_21 <= _GEN_103;
      end
    end else begin
      flight_21 <= _GEN_103;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_22 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h16 == auto_out_d_bits_source) begin
        flight_22 <= 1'h0;
      end else begin
        flight_22 <= _GEN_104;
      end
    end else begin
      flight_22 <= _GEN_104;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_23 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h17 == auto_out_d_bits_source) begin
        flight_23 <= 1'h0;
      end else begin
        flight_23 <= _GEN_105;
      end
    end else begin
      flight_23 <= _GEN_105;
    end
    if (_stalls_id_T_29) begin // @[Reg.scala 17:18]
      stalls_id_7 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_24 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h18 == auto_out_d_bits_source) begin
        flight_24 <= 1'h0;
      end else begin
        flight_24 <= _GEN_106;
      end
    end else begin
      flight_24 <= _GEN_106;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_25 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h19 == auto_out_d_bits_source) begin
        flight_25 <= 1'h0;
      end else begin
        flight_25 <= _GEN_107;
      end
    end else begin
      flight_25 <= _GEN_107;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_26 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h1a == auto_out_d_bits_source) begin
        flight_26 <= 1'h0;
      end else begin
        flight_26 <= _GEN_108;
      end
    end else begin
      flight_26 <= _GEN_108;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_27 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h1b == auto_out_d_bits_source) begin
        flight_27 <= 1'h0;
      end else begin
        flight_27 <= _GEN_109;
      end
    end else begin
      flight_27 <= _GEN_109;
    end
    if (_stalls_id_T_33) begin // @[Reg.scala 17:18]
      stalls_id_8 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_28 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h1c == auto_out_d_bits_source) begin
        flight_28 <= 1'h0;
      end else begin
        flight_28 <= _GEN_110;
      end
    end else begin
      flight_28 <= _GEN_110;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_29 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h1d == auto_out_d_bits_source) begin
        flight_29 <= 1'h0;
      end else begin
        flight_29 <= _GEN_111;
      end
    end else begin
      flight_29 <= _GEN_111;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_30 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h1e == auto_out_d_bits_source) begin
        flight_30 <= 1'h0;
      end else begin
        flight_30 <= _GEN_112;
      end
    end else begin
      flight_30 <= _GEN_112;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_31 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h1f == auto_out_d_bits_source) begin
        flight_31 <= 1'h0;
      end else begin
        flight_31 <= _GEN_113;
      end
    end else begin
      flight_31 <= _GEN_113;
    end
    if (_stalls_id_T_37) begin // @[Reg.scala 17:18]
      stalls_id_9 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_32 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h20 == auto_out_d_bits_source) begin
        flight_32 <= 1'h0;
      end else begin
        flight_32 <= _GEN_114;
      end
    end else begin
      flight_32 <= _GEN_114;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_33 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h21 == auto_out_d_bits_source) begin
        flight_33 <= 1'h0;
      end else begin
        flight_33 <= _GEN_115;
      end
    end else begin
      flight_33 <= _GEN_115;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_34 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h22 == auto_out_d_bits_source) begin
        flight_34 <= 1'h0;
      end else begin
        flight_34 <= _GEN_116;
      end
    end else begin
      flight_34 <= _GEN_116;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_35 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h23 == auto_out_d_bits_source) begin
        flight_35 <= 1'h0;
      end else begin
        flight_35 <= _GEN_117;
      end
    end else begin
      flight_35 <= _GEN_117;
    end
    if (_stalls_id_T_41) begin // @[Reg.scala 17:18]
      stalls_id_10 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_36 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h24 == auto_out_d_bits_source) begin
        flight_36 <= 1'h0;
      end else begin
        flight_36 <= _GEN_118;
      end
    end else begin
      flight_36 <= _GEN_118;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_37 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h25 == auto_out_d_bits_source) begin
        flight_37 <= 1'h0;
      end else begin
        flight_37 <= _GEN_119;
      end
    end else begin
      flight_37 <= _GEN_119;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_38 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h26 == auto_out_d_bits_source) begin
        flight_38 <= 1'h0;
      end else begin
        flight_38 <= _GEN_120;
      end
    end else begin
      flight_38 <= _GEN_120;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_39 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h27 == auto_out_d_bits_source) begin
        flight_39 <= 1'h0;
      end else begin
        flight_39 <= _GEN_121;
      end
    end else begin
      flight_39 <= _GEN_121;
    end
    if (_stalls_id_T_45) begin // @[Reg.scala 17:18]
      stalls_id_11 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_40 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h28 == auto_out_d_bits_source) begin
        flight_40 <= 1'h0;
      end else begin
        flight_40 <= _GEN_122;
      end
    end else begin
      flight_40 <= _GEN_122;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_41 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h29 == auto_out_d_bits_source) begin
        flight_41 <= 1'h0;
      end else begin
        flight_41 <= _GEN_123;
      end
    end else begin
      flight_41 <= _GEN_123;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_42 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h2a == auto_out_d_bits_source) begin
        flight_42 <= 1'h0;
      end else begin
        flight_42 <= _GEN_124;
      end
    end else begin
      flight_42 <= _GEN_124;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_43 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h2b == auto_out_d_bits_source) begin
        flight_43 <= 1'h0;
      end else begin
        flight_43 <= _GEN_125;
      end
    end else begin
      flight_43 <= _GEN_125;
    end
    if (_stalls_id_T_49) begin // @[Reg.scala 17:18]
      stalls_id_12 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_44 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h2c == auto_out_d_bits_source) begin
        flight_44 <= 1'h0;
      end else begin
        flight_44 <= _GEN_126;
      end
    end else begin
      flight_44 <= _GEN_126;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_45 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h2d == auto_out_d_bits_source) begin
        flight_45 <= 1'h0;
      end else begin
        flight_45 <= _GEN_127;
      end
    end else begin
      flight_45 <= _GEN_127;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_46 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h2e == auto_out_d_bits_source) begin
        flight_46 <= 1'h0;
      end else begin
        flight_46 <= _GEN_128;
      end
    end else begin
      flight_46 <= _GEN_128;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_47 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h2f == auto_out_d_bits_source) begin
        flight_47 <= 1'h0;
      end else begin
        flight_47 <= _GEN_129;
      end
    end else begin
      flight_47 <= _GEN_129;
    end
    if (_stalls_id_T_53) begin // @[Reg.scala 17:18]
      stalls_id_13 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_48 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h30 == auto_out_d_bits_source) begin
        flight_48 <= 1'h0;
      end else begin
        flight_48 <= _GEN_130;
      end
    end else begin
      flight_48 <= _GEN_130;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_49 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h31 == auto_out_d_bits_source) begin
        flight_49 <= 1'h0;
      end else begin
        flight_49 <= _GEN_131;
      end
    end else begin
      flight_49 <= _GEN_131;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_50 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h32 == auto_out_d_bits_source) begin
        flight_50 <= 1'h0;
      end else begin
        flight_50 <= _GEN_132;
      end
    end else begin
      flight_50 <= _GEN_132;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_51 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h33 == auto_out_d_bits_source) begin
        flight_51 <= 1'h0;
      end else begin
        flight_51 <= _GEN_133;
      end
    end else begin
      flight_51 <= _GEN_133;
    end
    if (_stalls_id_T_57) begin // @[Reg.scala 17:18]
      stalls_id_14 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_52 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h34 == auto_out_d_bits_source) begin
        flight_52 <= 1'h0;
      end else begin
        flight_52 <= _GEN_134;
      end
    end else begin
      flight_52 <= _GEN_134;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_53 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h35 == auto_out_d_bits_source) begin
        flight_53 <= 1'h0;
      end else begin
        flight_53 <= _GEN_135;
      end
    end else begin
      flight_53 <= _GEN_135;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_54 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h36 == auto_out_d_bits_source) begin
        flight_54 <= 1'h0;
      end else begin
        flight_54 <= _GEN_136;
      end
    end else begin
      flight_54 <= _GEN_136;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_55 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h37 == auto_out_d_bits_source) begin
        flight_55 <= 1'h0;
      end else begin
        flight_55 <= _GEN_137;
      end
    end else begin
      flight_55 <= _GEN_137;
    end
    if (_stalls_id_T_61) begin // @[Reg.scala 17:18]
      stalls_id_15 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_56 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h38 == auto_out_d_bits_source) begin
        flight_56 <= 1'h0;
      end else begin
        flight_56 <= _GEN_138;
      end
    end else begin
      flight_56 <= _GEN_138;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_57 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h39 == auto_out_d_bits_source) begin
        flight_57 <= 1'h0;
      end else begin
        flight_57 <= _GEN_139;
      end
    end else begin
      flight_57 <= _GEN_139;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_58 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h3a == auto_out_d_bits_source) begin
        flight_58 <= 1'h0;
      end else begin
        flight_58 <= _GEN_140;
      end
    end else begin
      flight_58 <= _GEN_140;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_59 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h3b == auto_out_d_bits_source) begin
        flight_59 <= 1'h0;
      end else begin
        flight_59 <= _GEN_141;
      end
    end else begin
      flight_59 <= _GEN_141;
    end
    if (_stalls_id_T_65) begin // @[Reg.scala 17:18]
      stalls_id_16 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_60 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h3c == auto_out_d_bits_source) begin
        flight_60 <= 1'h0;
      end else begin
        flight_60 <= _GEN_142;
      end
    end else begin
      flight_60 <= _GEN_142;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_61 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h3d == auto_out_d_bits_source) begin
        flight_61 <= 1'h0;
      end else begin
        flight_61 <= _GEN_143;
      end
    end else begin
      flight_61 <= _GEN_143;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_62 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h3e == auto_out_d_bits_source) begin
        flight_62 <= 1'h0;
      end else begin
        flight_62 <= _GEN_144;
      end
    end else begin
      flight_62 <= _GEN_144;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_63 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (7'h3f == auto_out_d_bits_source) begin
        flight_63 <= 1'h0;
      end else begin
        flight_63 <= _GEN_145;
      end
    end else begin
      flight_63 <= _GEN_145;
    end
    if (_stalls_id_T_69) begin // @[Reg.scala 17:18]
      stalls_id_17 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin
      if (d_first_first) begin
        if (d_first_beats1_opdata) begin
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    TLFIFOFixer_3_covState <= TLFIFOFixer_3_xor0;
    if (TLFIFOFixer_3_covMap_write_en & TLFIFOFixer_3_covMap_write_mask) begin
      TLFIFOFixer_3_covMap[TLFIFOFixer_3_covMap_write_addr] <= TLFIFOFixer_3_covMap_write_data; // @[Coverage map for TLFIFOFixer_3]
    end
    if (!(TLFIFOFixer_3_covMap_read_data | metaReset)) begin
      TLFIFOFixer_3_covSum <= TLFIFOFixer_3_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_101 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    TLFIFOFixer_3_covMap[initvar] = 0; //_101[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  flight_64 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  flight_65 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  flight_66 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  flight_67 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  flight_68 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  flight_69 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  flight_70 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  flight_71 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  stalls_id = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  flight_72 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  flight_73 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  flight_74 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  flight_75 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  flight_76 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  flight_77 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  flight_78 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  flight_79 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  stalls_id_1 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  flight_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  flight_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  flight_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  flight_3 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  stalls_id_2 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  flight_4 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  flight_5 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  flight_6 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  flight_7 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  stalls_id_3 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  flight_8 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  flight_9 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  flight_10 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  flight_11 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  stalls_id_4 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  flight_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  flight_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  flight_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  flight_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  stalls_id_5 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  flight_16 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  flight_17 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  flight_18 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  flight_19 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  stalls_id_6 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  flight_20 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  flight_21 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  flight_22 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  flight_23 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  stalls_id_7 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  flight_24 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  flight_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  flight_26 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  flight_27 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  stalls_id_8 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  flight_28 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  flight_29 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  flight_30 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  flight_31 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  stalls_id_9 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  flight_32 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  flight_33 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  flight_34 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  flight_35 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  stalls_id_10 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  flight_36 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  flight_37 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  flight_38 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  flight_39 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  stalls_id_11 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  flight_40 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  flight_41 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  flight_42 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  flight_43 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  stalls_id_12 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  flight_44 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  flight_45 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  flight_46 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  flight_47 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  stalls_id_13 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  flight_48 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  flight_49 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  flight_50 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  flight_51 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  stalls_id_14 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  flight_52 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  flight_53 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  flight_54 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  flight_55 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  stalls_id_15 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  flight_56 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  flight_57 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  flight_58 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  flight_59 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  stalls_id_16 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  flight_60 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  flight_61 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  flight_62 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  flight_63 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  stalls_id_17 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  d_first_counter = _RAND_99[8:0];
  _RAND_100 = {1{`RANDOM}};
  TLFIFOFixer_3_covState = 0; //_100[19:0];
  _RAND_102 = {1{`RANDOM}};
  TLFIFOFixer_3_covSum = 0; //_102[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar_5(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [30:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_6_a_ready,
  output        auto_out_6_a_valid,
  output [2:0]  auto_out_6_a_bits_opcode,
  output [2:0]  auto_out_6_a_bits_size,
  output [6:0]  auto_out_6_a_bits_source,
  output [11:0] auto_out_6_a_bits_address,
  output [7:0]  auto_out_6_a_bits_mask,
  output        auto_out_6_d_ready,
  input         auto_out_6_d_valid,
  input  [2:0]  auto_out_6_d_bits_opcode,
  input  [2:0]  auto_out_6_d_bits_size,
  input  [6:0]  auto_out_6_d_bits_source,
  input  [63:0] auto_out_6_d_bits_data,
  input         auto_out_5_a_ready,
  output        auto_out_5_a_valid,
  output [2:0]  auto_out_5_a_bits_size,
  output [6:0]  auto_out_5_a_bits_source,
  output [17:0] auto_out_5_a_bits_address,
  output [7:0]  auto_out_5_a_bits_mask,
  output        auto_out_5_d_ready,
  input         auto_out_5_d_valid,
  input  [2:0]  auto_out_5_d_bits_size,
  input  [6:0]  auto_out_5_d_bits_source,
  input  [63:0] auto_out_5_d_bits_data,
  input         auto_out_4_a_ready,
  output        auto_out_4_a_valid,
  output [2:0]  auto_out_4_a_bits_size,
  output [6:0]  auto_out_4_a_bits_source,
  output [16:0] auto_out_4_a_bits_address,
  output [7:0]  auto_out_4_a_bits_mask,
  output        auto_out_4_d_ready,
  input         auto_out_4_d_valid,
  input  [2:0]  auto_out_4_d_bits_size,
  input  [6:0]  auto_out_4_d_bits_source,
  input  [63:0] auto_out_4_d_bits_data,
  input         auto_out_3_a_ready,
  output        auto_out_3_a_valid,
  output [2:0]  auto_out_3_a_bits_opcode,
  output [2:0]  auto_out_3_a_bits_size,
  output [6:0]  auto_out_3_a_bits_source,
  output [25:0] auto_out_3_a_bits_address,
  output [7:0]  auto_out_3_a_bits_mask,
  output [63:0] auto_out_3_a_bits_data,
  output        auto_out_3_d_ready,
  input         auto_out_3_d_valid,
  input  [2:0]  auto_out_3_d_bits_opcode,
  input  [2:0]  auto_out_3_d_bits_size,
  input  [6:0]  auto_out_3_d_bits_source,
  input  [63:0] auto_out_3_d_bits_data,
  input         auto_out_2_a_ready,
  output        auto_out_2_a_valid,
  output [2:0]  auto_out_2_a_bits_opcode,
  output [2:0]  auto_out_2_a_bits_size,
  output [6:0]  auto_out_2_a_bits_source,
  output [27:0] auto_out_2_a_bits_address,
  output [7:0]  auto_out_2_a_bits_mask,
  output [63:0] auto_out_2_a_bits_data,
  output        auto_out_2_d_ready,
  input         auto_out_2_d_valid,
  input  [2:0]  auto_out_2_d_bits_opcode,
  input  [2:0]  auto_out_2_d_bits_size,
  input  [6:0]  auto_out_2_d_bits_source,
  input  [63:0] auto_out_2_d_bits_data,
  input         auto_out_1_a_ready,
  output        auto_out_1_a_valid,
  output [2:0]  auto_out_1_a_bits_opcode,
  output [2:0]  auto_out_1_a_bits_param,
  output [2:0]  auto_out_1_a_bits_size,
  output [6:0]  auto_out_1_a_bits_source,
  output [30:0] auto_out_1_a_bits_address,
  output [7:0]  auto_out_1_a_bits_mask,
  output [63:0] auto_out_1_a_bits_data,
  output        auto_out_1_d_ready,
  input         auto_out_1_d_valid,
  input  [2:0]  auto_out_1_d_bits_opcode,
  input  [2:0]  auto_out_1_d_bits_size,
  input  [6:0]  auto_out_1_d_bits_source,
  input         auto_out_1_d_bits_denied,
  input  [63:0] auto_out_1_d_bits_data,
  input         auto_out_1_d_bits_corrupt,
  input         auto_out_0_a_ready,
  output        auto_out_0_a_valid,
  output [2:0]  auto_out_0_a_bits_opcode,
  output [3:0]  auto_out_0_a_bits_size,
  output [6:0]  auto_out_0_a_bits_source,
  output        auto_out_0_d_ready,
  input         auto_out_0_d_valid,
  input  [2:0]  auto_out_0_d_bits_opcode,
  input  [3:0]  auto_out_0_d_bits_size,
  input  [6:0]  auto_out_0_d_bits_source,
  input         auto_out_0_d_bits_denied,
  input  [63:0] auto_out_0_d_bits_data,
  input         auto_out_0_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 9'h0; // @[Arbiter.scala 88:28]
  wire [6:0] readys_valid = {auto_out_6_d_valid,auto_out_5_d_valid,auto_out_4_d_valid,auto_out_3_d_valid,
    auto_out_2_d_valid,auto_out_1_d_valid,auto_out_0_d_valid}; // @[Cat.scala 31:58]
  reg [6:0] readys_mask; // @[Arbiter.scala 23:23]
  wire [6:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 24:30]
  wire [6:0] _readys_filter_T_1 = readys_valid & _readys_filter_T; // @[Arbiter.scala 24:28]
  wire [13:0] readys_filter = {_readys_filter_T_1,auto_out_6_d_valid,auto_out_5_d_valid,auto_out_4_d_valid,
    auto_out_3_d_valid,auto_out_2_d_valid,auto_out_1_d_valid,auto_out_0_d_valid}; // @[Cat.scala 31:58]
  wire [13:0] _GEN_1 = {{1'd0}, readys_filter[13:1]}; // @[package.scala 253:43]
  wire [13:0] _readys_unready_T_1 = readys_filter | _GEN_1; // @[package.scala 253:43]
  wire [13:0] _GEN_2 = {{2'd0}, _readys_unready_T_1[13:2]}; // @[package.scala 253:43]
  wire [13:0] _readys_unready_T_3 = _readys_unready_T_1 | _GEN_2; // @[package.scala 253:43]
  wire [13:0] _GEN_3 = {{4'd0}, _readys_unready_T_3[13:4]}; // @[package.scala 253:43]
  wire [13:0] _readys_unready_T_5 = _readys_unready_T_3 | _GEN_3; // @[package.scala 253:43]
  wire [13:0] _readys_unready_T_8 = {readys_mask, 7'h0}; // @[Arbiter.scala 25:66]
  wire [13:0] _GEN_4 = {{1'd0}, _readys_unready_T_5[13:1]}; // @[Arbiter.scala 25:58]
  wire [13:0] readys_unready = _GEN_4 | _readys_unready_T_8; // @[Arbiter.scala 25:58]
  wire [6:0] _readys_readys_T_2 = readys_unready[13:7] & readys_unready[6:0]; // @[Arbiter.scala 26:39]
  wire [6:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 26:18]
  wire  readys_0 = readys_readys[0]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_0 = readys_0 & auto_out_0_d_valid; // @[Arbiter.scala 97:79]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire [6:0] _T_116 = muxStateEarly_0 ? auto_out_0_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire  readys_1 = readys_readys[1]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_1 = readys_1 & auto_out_1_d_valid; // @[Arbiter.scala 97:79]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire [6:0] _T_117 = muxStateEarly_1 ? auto_out_1_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_123 = _T_116 | _T_117; // @[Mux.scala 27:73]
  wire  readys_2 = readys_readys[2]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_2 = readys_2 & auto_out_2_d_valid; // @[Arbiter.scala 97:79]
  reg  state_2; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_2 = idle ? earlyWinner_2 : state_2; // @[Arbiter.scala 117:30]
  wire [6:0] _T_118 = muxStateEarly_2 ? auto_out_2_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_124 = _T_123 | _T_118; // @[Mux.scala 27:73]
  wire  readys_3 = readys_readys[3]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_3 = readys_3 & auto_out_3_d_valid; // @[Arbiter.scala 97:79]
  reg  state_3; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_3 = idle ? earlyWinner_3 : state_3; // @[Arbiter.scala 117:30]
  wire [6:0] _T_119 = muxStateEarly_3 ? auto_out_3_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_125 = _T_124 | _T_119; // @[Mux.scala 27:73]
  wire  readys_4 = readys_readys[4]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_4 = readys_4 & auto_out_4_d_valid; // @[Arbiter.scala 97:79]
  reg  state_4; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_4 = idle ? earlyWinner_4 : state_4; // @[Arbiter.scala 117:30]
  wire [6:0] _T_120 = muxStateEarly_4 ? auto_out_4_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_126 = _T_125 | _T_120; // @[Mux.scala 27:73]
  wire  readys_5 = readys_readys[5]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_5 = readys_5 & auto_out_5_d_valid; // @[Arbiter.scala 97:79]
  reg  state_5; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_5 = idle ? earlyWinner_5 : state_5; // @[Arbiter.scala 117:30]
  wire [6:0] _T_121 = muxStateEarly_5 ? auto_out_5_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_127 = _T_126 | _T_121; // @[Mux.scala 27:73]
  wire  readys_6 = readys_readys[6]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_6 = readys_6 & auto_out_6_d_valid; // @[Arbiter.scala 97:79]
  reg  state_6; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_6 = idle ? earlyWinner_6 : state_6; // @[Arbiter.scala 117:30]
  wire [6:0] _T_122 = muxStateEarly_6 ? auto_out_6_d_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [30:0] _requestAIO_T = auto_in_a_bits_address ^ 31'h2000; // @[Parameters.scala 137:31]
  wire [31:0] _requestAIO_T_1 = {1'b0,$signed(_requestAIO_T)}; // @[Parameters.scala 137:49]
  wire [31:0] _requestAIO_T_3 = $signed(_requestAIO_T_1) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_0 = $signed(_requestAIO_T_3) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _requestAIO_T_5 = auto_in_a_bits_address ^ 31'h44000000; // @[Parameters.scala 137:31]
  wire [31:0] _requestAIO_T_6 = {1'b0,$signed(_requestAIO_T_5)}; // @[Parameters.scala 137:49]
  wire [31:0] _requestAIO_T_8 = $signed(_requestAIO_T_6) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_1 = $signed(_requestAIO_T_8) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _requestAIO_T_10 = auto_in_a_bits_address ^ 31'h4000000; // @[Parameters.scala 137:31]
  wire [31:0] _requestAIO_T_11 = {1'b0,$signed(_requestAIO_T_10)}; // @[Parameters.scala 137:49]
  wire [31:0] _requestAIO_T_13 = $signed(_requestAIO_T_11) & 32'sh44000000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_2 = $signed(_requestAIO_T_13) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _requestAIO_T_15 = auto_in_a_bits_address ^ 31'h2000000; // @[Parameters.scala 137:31]
  wire [31:0] _requestAIO_T_16 = {1'b0,$signed(_requestAIO_T_15)}; // @[Parameters.scala 137:49]
  wire [31:0] _requestAIO_T_18 = $signed(_requestAIO_T_16) & 32'sh46030000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_3 = $signed(_requestAIO_T_18) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _requestAIO_T_20 = auto_in_a_bits_address ^ 31'h10000; // @[Parameters.scala 137:31]
  wire [31:0] _requestAIO_T_21 = {1'b0,$signed(_requestAIO_T_20)}; // @[Parameters.scala 137:49]
  wire [31:0] _requestAIO_T_23 = $signed(_requestAIO_T_21) & 32'sh46030000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_4 = $signed(_requestAIO_T_23) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _requestAIO_T_25 = auto_in_a_bits_address ^ 31'h20000; // @[Parameters.scala 137:31]
  wire [31:0] _requestAIO_T_26 = {1'b0,$signed(_requestAIO_T_25)}; // @[Parameters.scala 137:49]
  wire [31:0] _requestAIO_T_28 = $signed(_requestAIO_T_26) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_5 = $signed(_requestAIO_T_28) == 32'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _requestAIO_T_31 = {1'b0,$signed(auto_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [31:0] _requestAIO_T_33 = $signed(_requestAIO_T_31) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  requestAIO_0_6 = $signed(_requestAIO_T_33) == 32'sh0; // @[Parameters.scala 137:67]
  wire [26:0] _beatsDO_decode_T_1 = 27'hfff << auto_out_0_d_bits_size; // @[package.scala 234:77]
  wire [11:0] _beatsDO_decode_T_3 = ~_beatsDO_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] beatsDO_decode = _beatsDO_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata = auto_out_0_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [8:0] beatsDO_0 = beatsDO_opdata ? beatsDO_decode : 9'h0; // @[Edges.scala 220:14]
  wire [3:0] out_1_1_d_bits_size = {{1'd0}, auto_out_1_d_bits_size}; // @[BundleMap.scala 247:19 Xbar.scala 288:19]
  wire [20:0] _beatsDO_decode_T_5 = 21'h3f << out_1_1_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_7 = ~_beatsDO_decode_T_5[5:0]; // @[package.scala 234:46]
  wire [2:0] beatsDO_decode_1 = _beatsDO_decode_T_7[5:3]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata_1 = auto_out_1_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] beatsDO_1 = beatsDO_opdata_1 ? beatsDO_decode_1 : 3'h0; // @[Edges.scala 220:14]
  wire [3:0] out_1_2_d_bits_size = {{1'd0}, auto_out_2_d_bits_size}; // @[BundleMap.scala 247:19 Xbar.scala 288:19]
  wire [20:0] _beatsDO_decode_T_9 = 21'h3f << out_1_2_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_11 = ~_beatsDO_decode_T_9[5:0]; // @[package.scala 234:46]
  wire [2:0] beatsDO_decode_2 = _beatsDO_decode_T_11[5:3]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata_2 = auto_out_2_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] beatsDO_2 = beatsDO_opdata_2 ? beatsDO_decode_2 : 3'h0; // @[Edges.scala 220:14]
  wire [3:0] out_1_3_d_bits_size = {{1'd0}, auto_out_3_d_bits_size}; // @[BundleMap.scala 247:19 Xbar.scala 288:19]
  wire [20:0] _beatsDO_decode_T_13 = 21'h3f << out_1_3_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_15 = ~_beatsDO_decode_T_13[5:0]; // @[package.scala 234:46]
  wire [2:0] beatsDO_decode_3 = _beatsDO_decode_T_15[5:3]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata_3 = auto_out_3_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] beatsDO_3 = beatsDO_opdata_3 ? beatsDO_decode_3 : 3'h0; // @[Edges.scala 220:14]
  wire [3:0] out_1_4_d_bits_size = {{1'd0}, auto_out_4_d_bits_size}; // @[BundleMap.scala 247:19 Xbar.scala 288:19]
  wire [20:0] _beatsDO_decode_T_17 = 21'h3f << out_1_4_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_19 = ~_beatsDO_decode_T_17[5:0]; // @[package.scala 234:46]
  wire [2:0] beatsDO_decode_4 = _beatsDO_decode_T_19[5:3]; // @[Edges.scala 219:59]
  wire [3:0] out_1_5_d_bits_size = {{1'd0}, auto_out_5_d_bits_size}; // @[BundleMap.scala 247:19 Xbar.scala 288:19]
  wire [20:0] _beatsDO_decode_T_21 = 21'h3f << out_1_5_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_23 = ~_beatsDO_decode_T_21[5:0]; // @[package.scala 234:46]
  wire [2:0] beatsDO_decode_5 = _beatsDO_decode_T_23[5:3]; // @[Edges.scala 219:59]
  wire [3:0] out_1_6_d_bits_size = {{1'd0}, auto_out_6_d_bits_size}; // @[BundleMap.scala 247:19 Xbar.scala 288:19]
  wire [20:0] _beatsDO_decode_T_25 = 21'h3f << out_1_6_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beatsDO_decode_T_27 = ~_beatsDO_decode_T_25[5:0]; // @[package.scala 234:46]
  wire [2:0] beatsDO_decode_6 = _beatsDO_decode_T_27[5:3]; // @[Edges.scala 219:59]
  wire  beatsDO_opdata_6 = auto_out_6_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] beatsDO_6 = beatsDO_opdata_6 ? beatsDO_decode_6 : 3'h0; // @[Edges.scala 220:14]
  wire  latch = idle & auto_in_d_ready; // @[Arbiter.scala 89:24]
  wire  _readys_T_3 = ~reset; // @[Arbiter.scala 22:12]
  wire [6:0] _readys_mask_T = readys_readys & readys_valid; // @[Arbiter.scala 28:29]
  wire [7:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 244:48]
  wire [6:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[6:0]; // @[package.scala 244:43]
  wire [8:0] _readys_mask_T_4 = {_readys_mask_T_3, 2'h0}; // @[package.scala 244:48]
  wire [6:0] _readys_mask_T_6 = _readys_mask_T_3 | _readys_mask_T_4[6:0]; // @[package.scala 244:43]
  wire [10:0] _readys_mask_T_7 = {_readys_mask_T_6, 4'h0}; // @[package.scala 244:48]
  wire [6:0] _readys_mask_T_9 = _readys_mask_T_6 | _readys_mask_T_7[6:0]; // @[package.scala 244:43]
  wire  prefixOR_2 = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 104:53]
  wire  prefixOR_3 = prefixOR_2 | earlyWinner_2; // @[Arbiter.scala 104:53]
  wire  prefixOR_4 = prefixOR_3 | earlyWinner_3; // @[Arbiter.scala 104:53]
  wire  prefixOR_5 = prefixOR_4 | earlyWinner_4; // @[Arbiter.scala 104:53]
  wire  prefixOR_6 = prefixOR_5 | earlyWinner_5; // @[Arbiter.scala 104:53]
  wire  _T_35 = auto_out_0_d_valid | auto_out_1_d_valid | auto_out_2_d_valid | auto_out_3_d_valid | auto_out_4_d_valid
     | auto_out_5_d_valid | auto_out_6_d_valid; // @[Arbiter.scala 107:36]
  wire  _T_36 = ~(auto_out_0_d_valid | auto_out_1_d_valid | auto_out_2_d_valid | auto_out_3_d_valid | auto_out_4_d_valid
     | auto_out_5_d_valid | auto_out_6_d_valid); // @[Arbiter.scala 107:15]
  wire [8:0] maskedBeats_0 = earlyWinner_0 ? beatsDO_0 : 9'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_1 = earlyWinner_1 ? beatsDO_1 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_2 = earlyWinner_2 ? beatsDO_2 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_3 = earlyWinner_3 ? beatsDO_3 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_4 = earlyWinner_4 ? beatsDO_decode_4 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_5 = earlyWinner_5 ? beatsDO_decode_5 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_6 = earlyWinner_6 ? beatsDO_6 : 3'h0; // @[Arbiter.scala 111:73]
  wire [8:0] _GEN_5 = {{6'd0}, maskedBeats_1}; // @[Arbiter.scala 112:44]
  wire [8:0] _initBeats_T = maskedBeats_0 | _GEN_5; // @[Arbiter.scala 112:44]
  wire [8:0] _GEN_6 = {{6'd0}, maskedBeats_2}; // @[Arbiter.scala 112:44]
  wire [8:0] _initBeats_T_1 = _initBeats_T | _GEN_6; // @[Arbiter.scala 112:44]
  wire [8:0] _GEN_7 = {{6'd0}, maskedBeats_3}; // @[Arbiter.scala 112:44]
  wire [8:0] _initBeats_T_2 = _initBeats_T_1 | _GEN_7; // @[Arbiter.scala 112:44]
  wire [8:0] _GEN_8 = {{6'd0}, maskedBeats_4}; // @[Arbiter.scala 112:44]
  wire [8:0] _initBeats_T_3 = _initBeats_T_2 | _GEN_8; // @[Arbiter.scala 112:44]
  wire [8:0] _GEN_9 = {{6'd0}, maskedBeats_5}; // @[Arbiter.scala 112:44]
  wire [8:0] _initBeats_T_4 = _initBeats_T_3 | _GEN_9; // @[Arbiter.scala 112:44]
  wire [8:0] _GEN_10 = {{6'd0}, maskedBeats_6}; // @[Arbiter.scala 112:44]
  wire [8:0] initBeats = _initBeats_T_4 | _GEN_10; // @[Arbiter.scala 112:44]
  wire  _sink_ACancel_earlyValid_T_18 = state_0 & auto_out_0_d_valid | state_1 & auto_out_1_d_valid | state_2 &
    auto_out_2_d_valid | state_3 & auto_out_3_d_valid | state_4 & auto_out_4_d_valid | state_5 & auto_out_5_d_valid |
    state_6 & auto_out_6_d_valid; // @[Mux.scala 27:73]
  wire  sink_ACancel_15_earlyValid = idle ? _T_35 : _sink_ACancel_earlyValid_T_18; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_15_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [8:0] _GEN_11 = {{8'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [8:0] _beatsLeft_T_4 = beatsLeft - _GEN_11; // @[Arbiter.scala 113:52]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  allowed_2 = idle ? readys_2 : state_2; // @[Arbiter.scala 121:24]
  wire  allowed_3 = idle ? readys_3 : state_3; // @[Arbiter.scala 121:24]
  wire  allowed_4 = idle ? readys_4 : state_4; // @[Arbiter.scala 121:24]
  wire  allowed_5 = idle ? readys_5 : state_5; // @[Arbiter.scala 121:24]
  wire  allowed_6 = idle ? readys_6 : state_6; // @[Arbiter.scala 121:24]
  wire [63:0] _T_77 = muxStateEarly_0 ? auto_out_0_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_78 = muxStateEarly_1 ? auto_out_1_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_79 = muxStateEarly_2 ? auto_out_2_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_80 = muxStateEarly_3 ? auto_out_3_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_81 = muxStateEarly_4 ? auto_out_4_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_82 = muxStateEarly_5 ? auto_out_5_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_83 = muxStateEarly_6 ? auto_out_6_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_84 = _T_77 | _T_78; // @[Mux.scala 27:73]
  wire [63:0] _T_85 = _T_84 | _T_79; // @[Mux.scala 27:73]
  wire [63:0] _T_86 = _T_85 | _T_80; // @[Mux.scala 27:73]
  wire [63:0] _T_87 = _T_86 | _T_81; // @[Mux.scala 27:73]
  wire [63:0] _T_88 = _T_87 | _T_82; // @[Mux.scala 27:73]
  wire [3:0] _T_129 = muxStateEarly_0 ? auto_out_0_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_130 = muxStateEarly_1 ? out_1_1_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_131 = muxStateEarly_2 ? out_1_2_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_132 = muxStateEarly_3 ? out_1_3_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_133 = muxStateEarly_4 ? out_1_4_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_134 = muxStateEarly_5 ? out_1_5_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_135 = muxStateEarly_6 ? out_1_6_d_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_136 = _T_129 | _T_130; // @[Mux.scala 27:73]
  wire [3:0] _T_137 = _T_136 | _T_131; // @[Mux.scala 27:73]
  wire [3:0] _T_138 = _T_137 | _T_132; // @[Mux.scala 27:73]
  wire [3:0] _T_139 = _T_138 | _T_133; // @[Mux.scala 27:73]
  wire [3:0] _T_140 = _T_139 | _T_134; // @[Mux.scala 27:73]
  wire [2:0] _T_155 = muxStateEarly_0 ? auto_out_0_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_156 = muxStateEarly_1 ? auto_out_1_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_157 = muxStateEarly_2 ? auto_out_2_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_158 = muxStateEarly_3 ? auto_out_3_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_159 = muxStateEarly_4 ? 3'h1 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_160 = muxStateEarly_5 ? 3'h1 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_161 = muxStateEarly_6 ? auto_out_6_d_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_162 = _T_155 | _T_156; // @[Mux.scala 27:73]
  wire [2:0] _T_163 = _T_162 | _T_157; // @[Mux.scala 27:73]
  wire [2:0] _T_164 = _T_163 | _T_158; // @[Mux.scala 27:73]
  wire [2:0] _T_165 = _T_164 | _T_159; // @[Mux.scala 27:73]
  wire [2:0] _T_166 = _T_165 | _T_160; // @[Mux.scala 27:73]
  reg  TLXbar_5_covState; // @[Register tracking TLXbar_5 state]
  reg  TLXbar_5_covMap [0:1]; // @[Coverage map for TLXbar_5]
  wire  TLXbar_5_covMap_read_en; // @[Coverage map for TLXbar_5]
  wire  TLXbar_5_covMap_read_addr; // @[Coverage map for TLXbar_5]
  wire  TLXbar_5_covMap_read_data; // @[Coverage map for TLXbar_5]
  wire  TLXbar_5_covMap_write_data; // @[Coverage map for TLXbar_5]
  wire  TLXbar_5_covMap_write_addr; // @[Coverage map for TLXbar_5]
  wire  TLXbar_5_covMap_write_mask; // @[Coverage map for TLXbar_5]
  wire  TLXbar_5_covMap_write_en; // @[Coverage map for TLXbar_5]
  reg [29:0] TLXbar_5_covSum; // @[Sum of coverage map]
  wire  state_2_shl;
  wire  state_2_pad;
  wire  state_3_shl;
  wire  state_3_pad;
  wire  state_4_shl;
  wire  state_4_pad;
  wire  state_5_shl;
  wire  state_5_pad;
  wire  state_1_shl;
  wire  state_1_pad;
  wire  state_0_shl;
  wire  state_0_pad;
  wire  state_6_shl;
  wire  state_6_pad;
  wire  TLXbar_5_xor4;
  wire  TLXbar_5_xor1;
  wire  TLXbar_5_xor5;
  wire  TLXbar_5_xor6;
  wire  TLXbar_5_xor2;
  wire  TLXbar_5_xor0;
  assign auto_in_a_ready = requestAIO_0_0 & auto_out_0_a_ready | requestAIO_0_1 & auto_out_1_a_ready | requestAIO_0_2 &
    auto_out_2_a_ready | requestAIO_0_3 & auto_out_3_a_ready | requestAIO_0_4 & auto_out_4_a_ready | requestAIO_0_5 &
    auto_out_5_a_ready | requestAIO_0_6 & auto_out_6_a_ready; // @[Mux.scala 27:73]
  assign auto_in_d_valid = idle ? _T_35 : _sink_ACancel_earlyValid_T_18; // @[Arbiter.scala 125:29]
  assign auto_in_d_bits_opcode = _T_166 | _T_161; // @[Mux.scala 27:73]
  assign auto_in_d_bits_size = _T_140 | _T_135; // @[Mux.scala 27:73]
  assign auto_in_d_bits_source = _T_127 | _T_122; // @[Mux.scala 27:73]
  assign auto_in_d_bits_denied = muxStateEarly_0 & auto_out_0_d_bits_denied | muxStateEarly_1 & auto_out_1_d_bits_denied
    ; // @[Mux.scala 27:73]
  assign auto_in_d_bits_data = _T_88 | _T_83; // @[Mux.scala 27:73]
  assign auto_in_d_bits_corrupt = muxStateEarly_0 & auto_out_0_d_bits_corrupt | muxStateEarly_1 &
    auto_out_1_d_bits_corrupt; // @[Mux.scala 27:73]
  assign auto_out_6_a_valid = auto_in_a_valid & requestAIO_0_6; // @[Xbar.scala 428:50]
  assign auto_out_6_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_6_a_bits_size = auto_in_a_bits_size[2:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_6_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_6_a_bits_address = auto_in_a_bits_address[11:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_6_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_6_d_ready = auto_in_d_ready & allowed_6; // @[Arbiter.scala 123:31]
  assign auto_out_5_a_valid = auto_in_a_valid & requestAIO_0_5; // @[Xbar.scala 428:50]
  assign auto_out_5_a_bits_size = auto_in_a_bits_size[2:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_5_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_5_a_bits_address = auto_in_a_bits_address[17:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_5_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_5_d_ready = auto_in_d_ready & allowed_5; // @[Arbiter.scala 123:31]
  assign auto_out_4_a_valid = auto_in_a_valid & requestAIO_0_4; // @[Xbar.scala 428:50]
  assign auto_out_4_a_bits_size = auto_in_a_bits_size[2:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_4_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_4_a_bits_address = auto_in_a_bits_address[16:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_4_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_4_d_ready = auto_in_d_ready & allowed_4; // @[Arbiter.scala 123:31]
  assign auto_out_3_a_valid = auto_in_a_valid & requestAIO_0_3; // @[Xbar.scala 428:50]
  assign auto_out_3_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_3_a_bits_size = auto_in_a_bits_size[2:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_3_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_3_a_bits_address = auto_in_a_bits_address[25:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_3_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_3_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_3_d_ready = auto_in_d_ready & allowed_3; // @[Arbiter.scala 123:31]
  assign auto_out_2_a_valid = auto_in_a_valid & requestAIO_0_2; // @[Xbar.scala 428:50]
  assign auto_out_2_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_2_a_bits_size = auto_in_a_bits_size[2:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_2_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_2_a_bits_address = auto_in_a_bits_address[27:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_2_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_2_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_2_d_ready = auto_in_d_ready & allowed_2; // @[Arbiter.scala 123:31]
  assign auto_out_1_a_valid = auto_in_a_valid & requestAIO_0_1; // @[Xbar.scala 428:50]
  assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_size = auto_in_a_bits_size[2:0]; // @[Xbar.scala 132:50 BundleMap.scala 247:19]
  assign auto_out_1_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_1_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1_d_ready = auto_in_d_ready & allowed_1; // @[Arbiter.scala 123:31]
  assign auto_out_0_a_valid = auto_in_a_valid & requestAIO_0_0; // @[Xbar.scala 428:50]
  assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_0_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign auto_out_0_d_ready = auto_in_d_ready & allowed_0; // @[Arbiter.scala 123:31]
  assign TLXbar_5_covMap_read_en = 1'h1;
  assign TLXbar_5_covMap_read_addr = TLXbar_5_covState;
  assign TLXbar_5_covMap_read_data = TLXbar_5_covMap[TLXbar_5_covMap_read_addr]; // @[Coverage map for TLXbar_5]
  assign TLXbar_5_covMap_write_data = 1'h1;
  assign TLXbar_5_covMap_write_addr = TLXbar_5_covState;
  assign TLXbar_5_covMap_write_mask = 1'h1;
  assign TLXbar_5_covMap_write_en = ~metaReset;
  assign state_2_shl = state_2;
  assign state_2_pad = state_2_shl;
  assign state_3_shl = state_3;
  assign state_3_pad = state_3_shl;
  assign state_4_shl = state_4;
  assign state_4_pad = state_4_shl;
  assign state_5_shl = state_5;
  assign state_5_pad = state_5_shl;
  assign state_1_shl = state_1;
  assign state_1_pad = state_1_shl;
  assign state_0_shl = state_0;
  assign state_0_pad = state_0_shl;
  assign state_6_shl = state_6;
  assign state_6_pad = state_6_shl;
  assign TLXbar_5_xor4 = state_3_pad ^ state_4_pad;
  assign TLXbar_5_xor1 = state_2_pad ^ TLXbar_5_xor4;
  assign TLXbar_5_xor5 = state_5_pad ^ state_1_pad;
  assign TLXbar_5_xor6 = state_0_pad ^ state_6_pad;
  assign TLXbar_5_xor2 = TLXbar_5_xor5 ^ TLXbar_5_xor6;
  assign TLXbar_5_xor0 = TLXbar_5_xor1 ^ TLXbar_5_xor2;
  assign io_covSum = TLXbar_5_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 9'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin
      beatsLeft <= initBeats;
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask <= 7'h7f; // @[Arbiter.scala 23:23]
    end else if (latch & |readys_valid) begin
      readys_mask <= _readys_mask_T_9;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_2 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_2 <= earlyWinner_2;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_3 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_3 <= earlyWinner_3;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_4 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_4 <= earlyWinner_4;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_5 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_5 <= earlyWinner_5;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_6 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_6 <= earlyWinner_6;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Arbiter.scala 22:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~((~earlyWinner_0 | ~earlyWinner_1) & (~prefixOR_2 | ~earlyWinner_2) & (~prefixOR_3 | ~earlyWinner_3) & (~
          prefixOR_4 | ~earlyWinner_4) & (~prefixOR_5 | ~earlyWinner_5) & (~prefixOR_6 | ~earlyWinner_6)) & _readys_T_3
          ) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~((~earlyWinner_0 | ~earlyWinner_1) & (~prefixOR_2 | ~earlyWinner_2) & (~prefixOR_3 | ~
          earlyWinner_3) & (~prefixOR_4 | ~earlyWinner_4) & (~prefixOR_5 | ~earlyWinner_5) & (~prefixOR_6 | ~
          earlyWinner_6))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(auto_out_0_d_valid | auto_out_1_d_valid | auto_out_2_d_valid | auto_out_3_d_valid | auto_out_4_d_valid
           | auto_out_5_d_valid | auto_out_6_d_valid) | (prefixOR_6 | earlyWinner_6)) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~(auto_out_0_d_valid | auto_out_1_d_valid | auto_out_2_d_valid | auto_out_3_d_valid |
          auto_out_4_d_valid | auto_out_5_d_valid | auto_out_6_d_valid) | (prefixOR_6 | earlyWinner_6))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_36 | _T_35) & _readys_T_3) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(_T_36 | _T_35)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    TLXbar_5_covState <= TLXbar_5_xor0;
    if (TLXbar_5_covMap_write_en & TLXbar_5_covMap_write_mask) begin
      TLXbar_5_covMap[TLXbar_5_covMap_write_addr] <= TLXbar_5_covMap_write_data; // @[Coverage map for TLXbar_5]
    end
    if (!(TLXbar_5_covMap_read_data | metaReset)) begin
      TLXbar_5_covSum <= TLXbar_5_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    TLXbar_5_covMap[initvar] = 0; //_10[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  readys_mask = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  state_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  TLXbar_5_covState = 0; //_9[0:0];
  _RAND_11 = {1{`RANDOM}};
  TLXbar_5_covSum = 0; //_11[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_13(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [30:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [30:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_param_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [6:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg [30:0] ram_address [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [30:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [30:0] ram_address_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_13_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_en = 1'h1;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_13_covSum = 30'h0;
  assign io_covSum = Queue_13_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= value_1 + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  value_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_14(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [3:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input         io_enq_bits_denied,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [3:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output        io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [6:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_denied [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_14_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_14_covSum = 30'h0;
  assign io_covSum = Queue_14_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= value_1 + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_5[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  value_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_4(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [30:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [30:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum
);
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_param; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire [30:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 361:21]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [30:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 361:21]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [29:0] bundleOut_0_a_q_io_covSum; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire [29:0] bundleIn_0_d_q_io_covSum; // @[Decoupled.scala 361:21]
  wire [29:0] TLBuffer_4_covSum;
  wire [29:0] bundleOut_0_a_q_sum;
  wire [29:0] bundleIn_0_d_q_sum;
  Queue_13 bundleOut_0_a_q ( // @[Decoupled.scala 361:21]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_covSum(bundleOut_0_a_q_io_covSum)
  );
  Queue_14 bundleIn_0_d_q ( // @[Decoupled.scala 361:21]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt),
    .io_covSum(bundleIn_0_d_q_io_covSum)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 Decoupled.scala 365:17]
  assign bundleOut_0_a_q_clock = clock;
  assign bundleOut_0_a_q_reset = reset;
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_clock = clock;
  assign bundleIn_0_d_q_reset = reset;
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBuffer_4_covSum = 30'h0;
  assign bundleOut_0_a_q_sum = TLBuffer_4_covSum + bundleOut_0_a_q_io_covSum;
  assign bundleIn_0_d_q_sum = bundleOut_0_a_q_sum + bundleIn_0_d_q_io_covSum;
  assign io_covSum = bundleIn_0_d_q_sum;
endmodule
module TLAtomicAutomata_1(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [30:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [30:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] cam_s_0_state; // @[AtomicAutomata.scala 76:28]
  reg [2:0] cam_a_0_bits_opcode; // @[AtomicAutomata.scala 77:24]
  reg [2:0] cam_a_0_bits_param; // @[AtomicAutomata.scala 77:24]
  reg [3:0] cam_a_0_bits_size; // @[AtomicAutomata.scala 77:24]
  reg [6:0] cam_a_0_bits_source; // @[AtomicAutomata.scala 77:24]
  reg [30:0] cam_a_0_bits_address; // @[AtomicAutomata.scala 77:24]
  reg [7:0] cam_a_0_bits_mask; // @[AtomicAutomata.scala 77:24]
  reg [63:0] cam_a_0_bits_data; // @[AtomicAutomata.scala 77:24]
  reg [3:0] cam_a_0_lut; // @[AtomicAutomata.scala 77:24]
  reg [63:0] cam_d_0_data; // @[AtomicAutomata.scala 78:24]
  reg  cam_d_0_denied; // @[AtomicAutomata.scala 78:24]
  reg  cam_d_0_corrupt; // @[AtomicAutomata.scala 78:24]
  wire  cam_free_0 = cam_s_0_state == 2'h0; // @[AtomicAutomata.scala 80:44]
  wire  cam_amo_0 = cam_s_0_state == 2'h2; // @[AtomicAutomata.scala 81:44]
  wire  cam_abusy_0 = cam_s_0_state == 2'h3 | cam_amo_0; // @[AtomicAutomata.scala 82:57]
  wire  cam_dmatch_0 = cam_s_0_state != 2'h0; // @[AtomicAutomata.scala 83:49]
  wire  _a_canLogical_T_1 = auto_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42]
  wire [30:0] _a_canLogical_T_4 = auto_in_a_bits_address ^ 31'h2000; // @[Parameters.scala 137:31]
  wire [31:0] _a_canLogical_T_5 = {1'b0,$signed(_a_canLogical_T_4)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_canLogical_T_7 = $signed(_a_canLogical_T_5) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  _a_canLogical_T_8 = $signed(_a_canLogical_T_7) == 32'sh0; // @[Parameters.scala 137:67]
  wire [30:0] _a_canLogical_T_9 = auto_in_a_bits_address ^ 31'h44000000; // @[Parameters.scala 137:31]
  wire [31:0] _a_canLogical_T_10 = {1'b0,$signed(_a_canLogical_T_9)}; // @[Parameters.scala 137:49]
  wire [31:0] _a_canLogical_T_12 = $signed(_a_canLogical_T_10) & 32'sh46032000; // @[Parameters.scala 137:52]
  wire  _a_canLogical_T_13 = $signed(_a_canLogical_T_12) == 32'sh0; // @[Parameters.scala 137:67]
  wire  _a_canLogical_T_14 = _a_canLogical_T_8 | _a_canLogical_T_13; // @[Parameters.scala 671:42]
  wire  a_canLogical = _a_canLogical_T_1 & _a_canLogical_T_14; // @[Parameters.scala 670:56]
  wire  a_isLogical = auto_in_a_bits_opcode == 3'h3; // @[AtomicAutomata.scala 90:47]
  wire  a_isArithmetic = auto_in_a_bits_opcode == 3'h2; // @[AtomicAutomata.scala 91:47]
  wire  _a_isSupported_T = a_isArithmetic ? a_canLogical : 1'h1; // @[AtomicAutomata.scala 92:63]
  wire  a_isSupported = a_isLogical ? a_canLogical : _a_isSupported_T; // @[AtomicAutomata.scala 92:32]
  wire [1:0] indexes_0 = {cam_a_0_bits_data[0],cam_d_0_data[0]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_1 = {cam_a_0_bits_data[1],cam_d_0_data[1]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_2 = {cam_a_0_bits_data[2],cam_d_0_data[2]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_3 = {cam_a_0_bits_data[3],cam_d_0_data[3]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_4 = {cam_a_0_bits_data[4],cam_d_0_data[4]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_5 = {cam_a_0_bits_data[5],cam_d_0_data[5]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_6 = {cam_a_0_bits_data[6],cam_d_0_data[6]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_7 = {cam_a_0_bits_data[7],cam_d_0_data[7]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_8 = {cam_a_0_bits_data[8],cam_d_0_data[8]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_9 = {cam_a_0_bits_data[9],cam_d_0_data[9]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_10 = {cam_a_0_bits_data[10],cam_d_0_data[10]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_11 = {cam_a_0_bits_data[11],cam_d_0_data[11]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_12 = {cam_a_0_bits_data[12],cam_d_0_data[12]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_13 = {cam_a_0_bits_data[13],cam_d_0_data[13]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_14 = {cam_a_0_bits_data[14],cam_d_0_data[14]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_15 = {cam_a_0_bits_data[15],cam_d_0_data[15]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_16 = {cam_a_0_bits_data[16],cam_d_0_data[16]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_17 = {cam_a_0_bits_data[17],cam_d_0_data[17]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_18 = {cam_a_0_bits_data[18],cam_d_0_data[18]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_19 = {cam_a_0_bits_data[19],cam_d_0_data[19]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_20 = {cam_a_0_bits_data[20],cam_d_0_data[20]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_21 = {cam_a_0_bits_data[21],cam_d_0_data[21]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_22 = {cam_a_0_bits_data[22],cam_d_0_data[22]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_23 = {cam_a_0_bits_data[23],cam_d_0_data[23]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_24 = {cam_a_0_bits_data[24],cam_d_0_data[24]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_25 = {cam_a_0_bits_data[25],cam_d_0_data[25]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_26 = {cam_a_0_bits_data[26],cam_d_0_data[26]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_27 = {cam_a_0_bits_data[27],cam_d_0_data[27]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_28 = {cam_a_0_bits_data[28],cam_d_0_data[28]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_29 = {cam_a_0_bits_data[29],cam_d_0_data[29]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_30 = {cam_a_0_bits_data[30],cam_d_0_data[30]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_31 = {cam_a_0_bits_data[31],cam_d_0_data[31]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_32 = {cam_a_0_bits_data[32],cam_d_0_data[32]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_33 = {cam_a_0_bits_data[33],cam_d_0_data[33]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_34 = {cam_a_0_bits_data[34],cam_d_0_data[34]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_35 = {cam_a_0_bits_data[35],cam_d_0_data[35]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_36 = {cam_a_0_bits_data[36],cam_d_0_data[36]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_37 = {cam_a_0_bits_data[37],cam_d_0_data[37]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_38 = {cam_a_0_bits_data[38],cam_d_0_data[38]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_39 = {cam_a_0_bits_data[39],cam_d_0_data[39]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_40 = {cam_a_0_bits_data[40],cam_d_0_data[40]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_41 = {cam_a_0_bits_data[41],cam_d_0_data[41]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_42 = {cam_a_0_bits_data[42],cam_d_0_data[42]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_43 = {cam_a_0_bits_data[43],cam_d_0_data[43]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_44 = {cam_a_0_bits_data[44],cam_d_0_data[44]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_45 = {cam_a_0_bits_data[45],cam_d_0_data[45]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_46 = {cam_a_0_bits_data[46],cam_d_0_data[46]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_47 = {cam_a_0_bits_data[47],cam_d_0_data[47]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_48 = {cam_a_0_bits_data[48],cam_d_0_data[48]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_49 = {cam_a_0_bits_data[49],cam_d_0_data[49]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_50 = {cam_a_0_bits_data[50],cam_d_0_data[50]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_51 = {cam_a_0_bits_data[51],cam_d_0_data[51]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_52 = {cam_a_0_bits_data[52],cam_d_0_data[52]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_53 = {cam_a_0_bits_data[53],cam_d_0_data[53]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_54 = {cam_a_0_bits_data[54],cam_d_0_data[54]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_55 = {cam_a_0_bits_data[55],cam_d_0_data[55]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_56 = {cam_a_0_bits_data[56],cam_d_0_data[56]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_57 = {cam_a_0_bits_data[57],cam_d_0_data[57]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_58 = {cam_a_0_bits_data[58],cam_d_0_data[58]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_59 = {cam_a_0_bits_data[59],cam_d_0_data[59]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_60 = {cam_a_0_bits_data[60],cam_d_0_data[60]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_61 = {cam_a_0_bits_data[61],cam_d_0_data[61]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_62 = {cam_a_0_bits_data[62],cam_d_0_data[62]}; // @[Cat.scala 31:58]
  wire [1:0] indexes_63 = {cam_a_0_bits_data[63],cam_d_0_data[63]}; // @[Cat.scala 31:58]
  wire [3:0] _logic_out_T = cam_a_0_lut >> indexes_0; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_2 = cam_a_0_lut >> indexes_1; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_4 = cam_a_0_lut >> indexes_2; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_6 = cam_a_0_lut >> indexes_3; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_8 = cam_a_0_lut >> indexes_4; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_10 = cam_a_0_lut >> indexes_5; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_12 = cam_a_0_lut >> indexes_6; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_14 = cam_a_0_lut >> indexes_7; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_16 = cam_a_0_lut >> indexes_8; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_18 = cam_a_0_lut >> indexes_9; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_20 = cam_a_0_lut >> indexes_10; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_22 = cam_a_0_lut >> indexes_11; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_24 = cam_a_0_lut >> indexes_12; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_26 = cam_a_0_lut >> indexes_13; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_28 = cam_a_0_lut >> indexes_14; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_30 = cam_a_0_lut >> indexes_15; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_32 = cam_a_0_lut >> indexes_16; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_34 = cam_a_0_lut >> indexes_17; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_36 = cam_a_0_lut >> indexes_18; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_38 = cam_a_0_lut >> indexes_19; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_40 = cam_a_0_lut >> indexes_20; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_42 = cam_a_0_lut >> indexes_21; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_44 = cam_a_0_lut >> indexes_22; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_46 = cam_a_0_lut >> indexes_23; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_48 = cam_a_0_lut >> indexes_24; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_50 = cam_a_0_lut >> indexes_25; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_52 = cam_a_0_lut >> indexes_26; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_54 = cam_a_0_lut >> indexes_27; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_56 = cam_a_0_lut >> indexes_28; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_58 = cam_a_0_lut >> indexes_29; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_60 = cam_a_0_lut >> indexes_30; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_62 = cam_a_0_lut >> indexes_31; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_64 = cam_a_0_lut >> indexes_32; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_66 = cam_a_0_lut >> indexes_33; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_68 = cam_a_0_lut >> indexes_34; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_70 = cam_a_0_lut >> indexes_35; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_72 = cam_a_0_lut >> indexes_36; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_74 = cam_a_0_lut >> indexes_37; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_76 = cam_a_0_lut >> indexes_38; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_78 = cam_a_0_lut >> indexes_39; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_80 = cam_a_0_lut >> indexes_40; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_82 = cam_a_0_lut >> indexes_41; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_84 = cam_a_0_lut >> indexes_42; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_86 = cam_a_0_lut >> indexes_43; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_88 = cam_a_0_lut >> indexes_44; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_90 = cam_a_0_lut >> indexes_45; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_92 = cam_a_0_lut >> indexes_46; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_94 = cam_a_0_lut >> indexes_47; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_96 = cam_a_0_lut >> indexes_48; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_98 = cam_a_0_lut >> indexes_49; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_100 = cam_a_0_lut >> indexes_50; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_102 = cam_a_0_lut >> indexes_51; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_104 = cam_a_0_lut >> indexes_52; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_106 = cam_a_0_lut >> indexes_53; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_108 = cam_a_0_lut >> indexes_54; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_110 = cam_a_0_lut >> indexes_55; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_112 = cam_a_0_lut >> indexes_56; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_114 = cam_a_0_lut >> indexes_57; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_116 = cam_a_0_lut >> indexes_58; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_118 = cam_a_0_lut >> indexes_59; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_120 = cam_a_0_lut >> indexes_60; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_122 = cam_a_0_lut >> indexes_61; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_124 = cam_a_0_lut >> indexes_62; // @[AtomicAutomata.scala 114:57]
  wire [3:0] _logic_out_T_126 = cam_a_0_lut >> indexes_63; // @[AtomicAutomata.scala 114:57]
  wire [7:0] logic_out_lo_lo_lo = {_logic_out_T_14[0],_logic_out_T_12[0],_logic_out_T_10[0],_logic_out_T_8[0],
    _logic_out_T_6[0],_logic_out_T_4[0],_logic_out_T_2[0],_logic_out_T[0]}; // @[Cat.scala 31:58]
  wire [15:0] logic_out_lo_lo = {_logic_out_T_30[0],_logic_out_T_28[0],_logic_out_T_26[0],_logic_out_T_24[0],
    _logic_out_T_22[0],_logic_out_T_20[0],_logic_out_T_18[0],_logic_out_T_16[0],logic_out_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] logic_out_lo_hi_lo = {_logic_out_T_46[0],_logic_out_T_44[0],_logic_out_T_42[0],_logic_out_T_40[0],
    _logic_out_T_38[0],_logic_out_T_36[0],_logic_out_T_34[0],_logic_out_T_32[0]}; // @[Cat.scala 31:58]
  wire [31:0] logic_out_lo = {_logic_out_T_62[0],_logic_out_T_60[0],_logic_out_T_58[0],_logic_out_T_56[0],
    _logic_out_T_54[0],_logic_out_T_52[0],_logic_out_T_50[0],_logic_out_T_48[0],logic_out_lo_hi_lo,logic_out_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] logic_out_hi_lo_lo = {_logic_out_T_78[0],_logic_out_T_76[0],_logic_out_T_74[0],_logic_out_T_72[0],
    _logic_out_T_70[0],_logic_out_T_68[0],_logic_out_T_66[0],_logic_out_T_64[0]}; // @[Cat.scala 31:58]
  wire [15:0] logic_out_hi_lo = {_logic_out_T_94[0],_logic_out_T_92[0],_logic_out_T_90[0],_logic_out_T_88[0],
    _logic_out_T_86[0],_logic_out_T_84[0],_logic_out_T_82[0],_logic_out_T_80[0],logic_out_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] logic_out_hi_hi_lo = {_logic_out_T_110[0],_logic_out_T_108[0],_logic_out_T_106[0],_logic_out_T_104[0],
    _logic_out_T_102[0],_logic_out_T_100[0],_logic_out_T_98[0],_logic_out_T_96[0]}; // @[Cat.scala 31:58]
  wire [31:0] logic_out_hi = {_logic_out_T_126[0],_logic_out_T_124[0],_logic_out_T_122[0],_logic_out_T_120[0],
    _logic_out_T_118[0],_logic_out_T_116[0],_logic_out_T_114[0],_logic_out_T_112[0],logic_out_hi_hi_lo,logic_out_hi_lo}; // @[Cat.scala 31:58]
  wire [63:0] logic_out = {logic_out_hi,logic_out_lo}; // @[Cat.scala 31:58]
  wire  unsigned_ = cam_a_0_bits_param[1]; // @[AtomicAutomata.scala 117:42]
  wire  take_max = cam_a_0_bits_param[0]; // @[AtomicAutomata.scala 118:42]
  wire  adder = cam_a_0_bits_param[2]; // @[AtomicAutomata.scala 119:39]
  wire [7:0] _signSel_T = ~cam_a_0_bits_mask; // @[AtomicAutomata.scala 121:25]
  wire [7:0] _GEN_10 = {{1'd0}, cam_a_0_bits_mask[7:1]}; // @[AtomicAutomata.scala 121:31]
  wire [7:0] _signSel_T_2 = _signSel_T | _GEN_10; // @[AtomicAutomata.scala 121:31]
  wire [7:0] signSel = ~_signSel_T_2; // @[AtomicAutomata.scala 121:23]
  wire [7:0] signbits_a = {cam_a_0_bits_data[63],cam_a_0_bits_data[55],cam_a_0_bits_data[47],cam_a_0_bits_data[39],
    cam_a_0_bits_data[31],cam_a_0_bits_data[23],cam_a_0_bits_data[15],cam_a_0_bits_data[7]}; // @[Cat.scala 31:58]
  wire [7:0] signbits_d = {cam_d_0_data[63],cam_d_0_data[55],cam_d_0_data[47],cam_d_0_data[39],cam_d_0_data[31],
    cam_d_0_data[23],cam_d_0_data[15],cam_d_0_data[7]}; // @[Cat.scala 31:58]
  wire [7:0] _signbit_a_T = signbits_a & signSel; // @[AtomicAutomata.scala 125:38]
  wire [8:0] _signbit_a_T_1 = {_signbit_a_T, 1'h0}; // @[AtomicAutomata.scala 125:49]
  wire [7:0] signbit_a = _signbit_a_T_1[7:0]; // @[AtomicAutomata.scala 125:54]
  wire [7:0] _signbit_d_T = signbits_d & signSel; // @[AtomicAutomata.scala 126:38]
  wire [8:0] _signbit_d_T_1 = {_signbit_d_T, 1'h0}; // @[AtomicAutomata.scala 126:49]
  wire [7:0] signbit_d = _signbit_d_T_1[7:0]; // @[AtomicAutomata.scala 126:54]
  wire [8:0] _signext_a_T = {signbit_a, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_a_T_2 = signbit_a | _signext_a_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _signext_a_T_3 = {_signext_a_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_a_T_5 = _signext_a_T_2 | _signext_a_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _signext_a_T_6 = {_signext_a_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_a_T_8 = _signext_a_T_5 | _signext_a_T_6[7:0]; // @[package.scala 244:43]
  wire [7:0] _signext_a_T_19 = _signext_a_T_8[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_21 = _signext_a_T_8[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_23 = _signext_a_T_8[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_25 = _signext_a_T_8[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_27 = _signext_a_T_8[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_29 = _signext_a_T_8[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_31 = _signext_a_T_8[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_a_T_33 = _signext_a_T_8[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] signext_a = {_signext_a_T_33,_signext_a_T_31,_signext_a_T_29,_signext_a_T_27,_signext_a_T_25,
    _signext_a_T_23,_signext_a_T_21,_signext_a_T_19}; // @[Cat.scala 31:58]
  wire [8:0] _signext_d_T = {signbit_d, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_d_T_2 = signbit_d | _signext_d_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _signext_d_T_3 = {_signext_d_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_d_T_5 = _signext_d_T_2 | _signext_d_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _signext_d_T_6 = {_signext_d_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _signext_d_T_8 = _signext_d_T_5 | _signext_d_T_6[7:0]; // @[package.scala 244:43]
  wire [7:0] _signext_d_T_19 = _signext_d_T_8[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_21 = _signext_d_T_8[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_23 = _signext_d_T_8[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_25 = _signext_d_T_8[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_27 = _signext_d_T_8[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_29 = _signext_d_T_8[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_31 = _signext_d_T_8[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _signext_d_T_33 = _signext_d_T_8[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] signext_d = {_signext_d_T_33,_signext_d_T_31,_signext_d_T_29,_signext_d_T_27,_signext_d_T_25,
    _signext_d_T_23,_signext_d_T_21,_signext_d_T_19}; // @[Cat.scala 31:58]
  wire [7:0] _wide_mask_T_9 = cam_a_0_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_11 = cam_a_0_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_13 = cam_a_0_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_15 = cam_a_0_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_17 = cam_a_0_bits_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_19 = cam_a_0_bits_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_21 = cam_a_0_bits_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _wide_mask_T_23 = cam_a_0_bits_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] wide_mask = {_wide_mask_T_23,_wide_mask_T_21,_wide_mask_T_19,_wide_mask_T_17,_wide_mask_T_15,
    _wide_mask_T_13,_wide_mask_T_11,_wide_mask_T_9}; // @[Cat.scala 31:58]
  wire [63:0] _a_a_ext_T = cam_a_0_bits_data & wide_mask; // @[AtomicAutomata.scala 131:28]
  wire [63:0] a_a_ext = _a_a_ext_T | signext_a; // @[AtomicAutomata.scala 131:41]
  wire [63:0] _a_d_ext_T = cam_d_0_data & wide_mask; // @[AtomicAutomata.scala 132:28]
  wire [63:0] a_d_ext = _a_d_ext_T | signext_d; // @[AtomicAutomata.scala 132:41]
  wire [63:0] _a_d_inv_T = ~a_d_ext; // @[AtomicAutomata.scala 133:43]
  wire [63:0] a_d_inv = adder ? a_d_ext : _a_d_inv_T; // @[AtomicAutomata.scala 133:26]
  wire [63:0] adder_out = a_a_ext + a_d_inv; // @[AtomicAutomata.scala 134:33]
  wire  a_bigger_uneq = unsigned_ == a_a_ext[63]; // @[AtomicAutomata.scala 136:38]
  wire  a_bigger = a_a_ext[63] == a_d_ext[63] ? ~adder_out[63] : a_bigger_uneq; // @[AtomicAutomata.scala 137:27]
  wire  pick_a = take_max == a_bigger; // @[AtomicAutomata.scala 138:31]
  wire [63:0] _arith_out_T = pick_a ? cam_a_0_bits_data : cam_d_0_data; // @[AtomicAutomata.scala 139:50]
  wire [63:0] arith_out = adder ? adder_out : _arith_out_T; // @[AtomicAutomata.scala 139:28]
  wire [63:0] amo_data = cam_a_0_bits_opcode[0] ? logic_out : arith_out; // @[AtomicAutomata.scala 145:14]
  wire  a_allow = ~cam_abusy_0 & (a_isSupported | cam_free_0); // @[AtomicAutomata.scala 149:35]
  reg [8:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 9'h0; // @[Arbiter.scala 88:28]
  wire  source_i_valid = auto_in_a_valid & a_allow; // @[AtomicAutomata.scala 151:38]
  wire [1:0] _readys_T = {source_i_valid,cam_amo_0}; // @[Cat.scala 31:58]
  wire [2:0] _readys_T_1 = {_readys_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0]; // @[package.scala 244:43]
  wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0}; // @[Arbiter.scala 16:78]
  wire [1:0] _readys_T_7 = ~_readys_T_5[1:0]; // @[Arbiter.scala 16:61]
  wire  readys_1 = _readys_T_7[1]; // @[Arbiter.scala 95:86]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 123:31]
  wire  _T = ~a_isSupported; // @[AtomicAutomata.scala 153:15]
  wire [2:0] source_i_bits_opcode = ~a_isSupported ? 3'h4 : auto_in_a_bits_opcode; // @[AtomicAutomata.scala 152:24 153:31 154:32]
  wire [2:0] source_i_bits_param = ~a_isSupported ? 3'h0 : auto_in_a_bits_param; // @[AtomicAutomata.scala 152:24 153:31 155:32]
  wire [1:0] source_c_bits_a_mask_sizeOH_shiftAmount = cam_a_0_bits_size[1:0]; // @[OneHot.scala 63:49]
  wire [3:0] _source_c_bits_a_mask_sizeOH_T_1 = 4'h1 << source_c_bits_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [2:0] source_c_bits_a_mask_sizeOH = _source_c_bits_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _source_c_bits_a_mask_T = cam_a_0_bits_size >= 4'h3; // @[Misc.scala 205:21]
  wire  source_c_bits_a_mask_size = source_c_bits_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  source_c_bits_a_mask_bit = cam_a_0_bits_address[2]; // @[Misc.scala 209:26]
  wire  source_c_bits_a_mask_nbit = ~source_c_bits_a_mask_bit; // @[Misc.scala 210:20]
  wire  source_c_bits_a_mask_acc = _source_c_bits_a_mask_T | source_c_bits_a_mask_size & source_c_bits_a_mask_nbit; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_acc_1 = _source_c_bits_a_mask_T | source_c_bits_a_mask_size & source_c_bits_a_mask_bit; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_size_1 = source_c_bits_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  source_c_bits_a_mask_bit_1 = cam_a_0_bits_address[1]; // @[Misc.scala 209:26]
  wire  source_c_bits_a_mask_nbit_1 = ~source_c_bits_a_mask_bit_1; // @[Misc.scala 210:20]
  wire  source_c_bits_a_mask_eq_2 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_2 = source_c_bits_a_mask_acc | source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_2; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_3 = source_c_bits_a_mask_nbit & source_c_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_3 = source_c_bits_a_mask_acc | source_c_bits_a_mask_size_1 & source_c_bits_a_mask_eq_3; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_4 = source_c_bits_a_mask_bit & source_c_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_4 = source_c_bits_a_mask_acc_1 | source_c_bits_a_mask_size_1 &
    source_c_bits_a_mask_eq_4; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_5 = source_c_bits_a_mask_bit & source_c_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_5 = source_c_bits_a_mask_acc_1 | source_c_bits_a_mask_size_1 &
    source_c_bits_a_mask_eq_5; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_size_2 = source_c_bits_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  source_c_bits_a_mask_bit_2 = cam_a_0_bits_address[0]; // @[Misc.scala 209:26]
  wire  source_c_bits_a_mask_nbit_2 = ~source_c_bits_a_mask_bit_2; // @[Misc.scala 210:20]
  wire  source_c_bits_a_mask_eq_6 = source_c_bits_a_mask_eq_2 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_6 = source_c_bits_a_mask_acc_2 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_6; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_7 = source_c_bits_a_mask_eq_2 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_7 = source_c_bits_a_mask_acc_2 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_7; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_8 = source_c_bits_a_mask_eq_3 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_8 = source_c_bits_a_mask_acc_3 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_8; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_9 = source_c_bits_a_mask_eq_3 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_9 = source_c_bits_a_mask_acc_3 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_9; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_10 = source_c_bits_a_mask_eq_4 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_10 = source_c_bits_a_mask_acc_4 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_10; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_11 = source_c_bits_a_mask_eq_4 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_11 = source_c_bits_a_mask_acc_4 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_11; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_12 = source_c_bits_a_mask_eq_5 & source_c_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_12 = source_c_bits_a_mask_acc_5 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_12; // @[Misc.scala 214:29]
  wire  source_c_bits_a_mask_eq_13 = source_c_bits_a_mask_eq_5 & source_c_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  source_c_bits_a_mask_acc_13 = source_c_bits_a_mask_acc_5 | source_c_bits_a_mask_size_2 &
    source_c_bits_a_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] source_c_bits_a_mask = {source_c_bits_a_mask_acc_13,source_c_bits_a_mask_acc_12,source_c_bits_a_mask_acc_11
    ,source_c_bits_a_mask_acc_10,source_c_bits_a_mask_acc_9,source_c_bits_a_mask_acc_8,source_c_bits_a_mask_acc_7,
    source_c_bits_a_mask_acc_6}; // @[Cat.scala 31:58]
  wire [26:0] _decode_T_1 = 27'hfff << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [11:0] _decode_T_3 = ~_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] decode = _decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 89:24]
  wire  readys_0 = _readys_T_7[0]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_0 = readys_0 & cam_amo_0; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1 = readys_1 & source_i_valid; // @[Arbiter.scala 97:79]
  wire  _T_10 = ~reset; // @[Arbiter.scala 105:13]
  wire  _T_12 = cam_amo_0 | source_i_valid; // @[Arbiter.scala 107:36]
  wire  _T_13 = ~(cam_amo_0 | source_i_valid); // @[Arbiter.scala 107:15]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & cam_amo_0 | state_1 & source_i_valid; // @[Mux.scala 27:73]
  wire  sink_ACancel_earlyValid = idle ? _T_12 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [8:0] _GEN_21 = {{8'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [8:0] _beatsLeft_T_4 = beatsLeft - _GEN_21; // @[Arbiter.scala 113:52]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  out_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 123:31]
  wire [63:0] _T_29 = muxStateEarly_0 ? amo_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_30 = muxStateEarly_1 ? auto_in_a_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_32 = muxStateEarly_0 ? source_c_bits_a_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_33 = muxStateEarly_1 ? auto_in_a_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [30:0] _T_35 = muxStateEarly_0 ? cam_a_0_bits_address : 31'h0; // @[Mux.scala 27:73]
  wire [30:0] _T_36 = muxStateEarly_1 ? auto_in_a_bits_address : 31'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_38 = muxStateEarly_0 ? cam_a_0_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _T_39 = muxStateEarly_1 ? auto_in_a_bits_source : 7'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_41 = muxStateEarly_0 ? cam_a_0_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_42 = muxStateEarly_1 ? auto_in_a_bits_size : 4'h0; // @[Mux.scala 27:73]
  wire  _T_50 = out_1_ready & source_i_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_39 = {{1'd0}, auto_in_a_bits_param[1:0]}; // @[Mux.scala 81:61]
  wire [3:0] _cam_a_0_lut_T_2 = 3'h1 == _GEN_39 ? 4'he : 4'h8; // @[Mux.scala 81:58]
  wire [1:0] _GEN_12 = cam_free_0 ? 2'h3 : cam_s_0_state; // @[AtomicAutomata.scala 187:23 188:23 76:28]
  wire [1:0] _GEN_23 = _T_50 & _T ? _GEN_12 : cam_s_0_state; // @[AtomicAutomata.scala 174:50 76:28]
  wire  _T_53 = out_ready & cam_amo_0; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_24 = cam_amo_0 ? 2'h1 : _GEN_23; // @[AtomicAutomata.scala 196:23 197:23]
  wire [1:0] _GEN_25 = _T_53 ? _GEN_24 : _GEN_23; // @[AtomicAutomata.scala 194:32]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27]
  wire  d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25]
  wire  d_ackd = auto_out_d_bits_opcode == 3'h1; // @[AtomicAutomata.scala 213:40]
  wire  d_cam_sel_raw_0 = cam_a_0_bits_source == auto_out_d_bits_source; // @[AtomicAutomata.scala 204:53]
  wire  d_cam_sel_match_0 = d_cam_sel_raw_0 & cam_dmatch_0; // @[AtomicAutomata.scala 205:83]
  wire  d_drop = d_first & d_ackd & d_cam_sel_match_0; // @[AtomicAutomata.scala 232:40]
  wire  bundleOut_0_d_ready = auto_in_d_ready | d_drop; // @[AtomicAutomata.scala 236:35]
  wire  _d_first_T = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28]
  wire  d_ack = auto_out_d_bits_opcode == 3'h0; // @[AtomicAutomata.scala 214:40]
  wire  d_replace = d_first & d_ack & d_cam_sel_match_0; // @[AtomicAutomata.scala 233:42]
  reg [2:0] TLAtomicAutomata_1_covState; // @[Register tracking TLAtomicAutomata_1 state]
  reg  TLAtomicAutomata_1_covMap [0:7]; // @[Coverage map for TLAtomicAutomata_1]
  wire  TLAtomicAutomata_1_covMap_read_en; // @[Coverage map for TLAtomicAutomata_1]
  wire [2:0] TLAtomicAutomata_1_covMap_read_addr; // @[Coverage map for TLAtomicAutomata_1]
  wire  TLAtomicAutomata_1_covMap_read_data; // @[Coverage map for TLAtomicAutomata_1]
  wire  TLAtomicAutomata_1_covMap_write_data; // @[Coverage map for TLAtomicAutomata_1]
  wire [2:0] TLAtomicAutomata_1_covMap_write_addr; // @[Coverage map for TLAtomicAutomata_1]
  wire  TLAtomicAutomata_1_covMap_write_mask; // @[Coverage map for TLAtomicAutomata_1]
  wire  TLAtomicAutomata_1_covMap_write_en; // @[Coverage map for TLAtomicAutomata_1]
  reg [29:0] TLAtomicAutomata_1_covSum; // @[Sum of coverage map]
  wire [1:0] cam_s_0_state_shl;
  wire [2:0] cam_s_0_state_pad;
  wire [2:0] state_0_shl;
  wire [2:0] state_0_pad;
  wire [2:0] state_1_shl;
  wire [2:0] state_1_pad;
  wire [2:0] TLAtomicAutomata_1_xor2;
  wire [2:0] TLAtomicAutomata_1_xor0;
  assign auto_in_a_ready = out_1_ready & a_allow; // @[AtomicAutomata.scala 150:38]
  assign auto_in_d_valid = auto_out_d_valid & ~d_drop; // @[AtomicAutomata.scala 235:35]
  assign auto_in_d_bits_opcode = d_replace ? 3'h1 : auto_out_d_bits_opcode; // @[AtomicAutomata.scala 238:19 239:26 240:28]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = d_replace ? cam_d_0_denied | auto_out_d_bits_denied : auto_out_d_bits_denied; // @[AtomicAutomata.scala 238:19 239:26 243:29]
  assign auto_in_d_bits_data = d_replace ? cam_d_0_data : auto_out_d_bits_data; // @[AtomicAutomata.scala 238:19 239:26 241:26]
  assign auto_in_d_bits_corrupt = d_replace ? cam_d_0_corrupt | auto_out_d_bits_denied : auto_out_d_bits_corrupt; // @[AtomicAutomata.scala 238:19 239:26 242:29]
  assign auto_out_a_valid = idle ? _T_12 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_out_a_bits_opcode = muxStateEarly_1 ? source_i_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  assign auto_out_a_bits_param = muxStateEarly_1 ? source_i_bits_param : 3'h0; // @[Mux.scala 27:73]
  assign auto_out_a_bits_size = _T_41 | _T_42; // @[Mux.scala 27:73]
  assign auto_out_a_bits_source = _T_38 | _T_39; // @[Mux.scala 27:73]
  assign auto_out_a_bits_address = _T_35 | _T_36; // @[Mux.scala 27:73]
  assign auto_out_a_bits_mask = _T_32 | _T_33; // @[Mux.scala 27:73]
  assign auto_out_a_bits_data = _T_29 | _T_30; // @[Mux.scala 27:73]
  assign auto_out_d_ready = auto_in_d_ready | d_drop; // @[AtomicAutomata.scala 236:35]
  assign TLAtomicAutomata_1_covMap_read_en = 1'h1;
  assign TLAtomicAutomata_1_covMap_read_addr = TLAtomicAutomata_1_covState;
  assign TLAtomicAutomata_1_covMap_read_data = TLAtomicAutomata_1_covMap[TLAtomicAutomata_1_covMap_read_addr]; // @[Coverage map for TLAtomicAutomata_1]
  assign TLAtomicAutomata_1_covMap_write_data = 1'h1;
  assign TLAtomicAutomata_1_covMap_write_addr = TLAtomicAutomata_1_covState;
  assign TLAtomicAutomata_1_covMap_write_mask = 1'h1;
  assign TLAtomicAutomata_1_covMap_write_en = ~metaReset;
  assign cam_s_0_state_shl = cam_s_0_state;
  assign cam_s_0_state_pad = {1'h0,cam_s_0_state_shl};
  assign state_0_shl = {state_0, 2'h0};
  assign state_0_pad = state_0_shl;
  assign state_1_shl = {state_1, 2'h0};
  assign state_1_pad = state_1_shl;
  assign TLAtomicAutomata_1_xor2 = state_0_pad ^ state_1_pad;
  assign TLAtomicAutomata_1_xor0 = cam_s_0_state_pad ^ TLAtomicAutomata_1_xor2;
  assign io_covSum = TLAtomicAutomata_1_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[AtomicAutomata.scala 76:28]
      cam_s_0_state <= 2'h0; // @[AtomicAutomata.scala 76:28]
    end else if (_d_first_T & d_first) begin
      if (d_cam_sel_match_0) begin
        if (d_ackd) begin
          cam_s_0_state <= 2'h2;
        end else begin
          cam_s_0_state <= 2'h0;
        end
      end else begin
        cam_s_0_state <= _GEN_25;
      end
    end else begin
      cam_s_0_state <= _GEN_25;
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_opcode <= auto_in_a_bits_opcode;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_param <= auto_in_a_bits_param;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_size <= auto_in_a_bits_size;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_source <= auto_in_a_bits_source;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_address <= auto_in_a_bits_address;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_mask <= auto_in_a_bits_mask;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        cam_a_0_bits_data <= auto_in_a_bits_data;
      end
    end
    if (_T_50 & _T) begin // @[AtomicAutomata.scala 174:50]
      if (cam_free_0) begin
        if (3'h3 == _GEN_39) begin
          cam_a_0_lut <= 4'hc;
        end else if (3'h0 == _GEN_39) begin
          cam_a_0_lut <= 4'h6;
        end else begin
          cam_a_0_lut <= _cam_a_0_lut_T_2;
        end
      end
    end
    if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0 & d_ackd) begin
        cam_d_0_data <= auto_out_d_bits_data;
      end
    end
    if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0 & d_ackd) begin
        cam_d_0_denied <= auto_out_d_bits_denied;
      end
    end
    if (_d_first_T & d_first) begin // @[AtomicAutomata.scala 216:40]
      if (d_cam_sel_match_0 & d_ackd) begin
        cam_d_0_corrupt <= auto_out_d_bits_corrupt;
      end
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 9'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin
      if (earlyWinner_1) begin
        if (opdata) begin
          beatsLeft <= decode;
        end else begin
          beatsLeft <= 9'h0;
        end
      end else begin
        beatsLeft <= 9'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin
      if (d_first) begin
        if (d_first_beats1_opdata) begin
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1) & ~reset) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~earlyWinner_0 | ~earlyWinner_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(cam_amo_0 | source_i_valid) | (earlyWinner_0 | earlyWinner_1)) & _T_10) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~(cam_amo_0 | source_i_valid) | (earlyWinner_0 | earlyWinner_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_13 | _T_12) & _T_10) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(_T_13 | _T_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    TLAtomicAutomata_1_covState <= TLAtomicAutomata_1_xor0;
    if (TLAtomicAutomata_1_covMap_write_en & TLAtomicAutomata_1_covMap_write_mask) begin
      TLAtomicAutomata_1_covMap[TLAtomicAutomata_1_covMap_write_addr] <= TLAtomicAutomata_1_covMap_write_data; // @[Coverage map for TLAtomicAutomata_1]
    end
    if (!(TLAtomicAutomata_1_covMap_read_data | metaReset)) begin
      TLAtomicAutomata_1_covSum <= TLAtomicAutomata_1_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    TLAtomicAutomata_1_covMap[initvar] = 0; //_17[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cam_s_0_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cam_a_0_bits_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  cam_a_0_bits_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  cam_a_0_bits_size = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  cam_a_0_bits_source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  cam_a_0_bits_address = _RAND_5[30:0];
  _RAND_6 = {1{`RANDOM}};
  cam_a_0_bits_mask = _RAND_6[7:0];
  _RAND_7 = {2{`RANDOM}};
  cam_a_0_bits_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  cam_a_0_lut = _RAND_8[3:0];
  _RAND_9 = {2{`RANDOM}};
  cam_d_0_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  cam_d_0_denied = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cam_d_0_corrupt = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  beatsLeft = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  state_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  d_first_counter = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  TLAtomicAutomata_1_covState = 0; //_16[2:0];
  _RAND_18 = {1{`RANDOM}};
  TLAtomicAutomata_1_covSum = 0; //_18[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_15(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [3:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [3:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [6:0] ram_source [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_15_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = 1'h0;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = 1'h0;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_15_covSum = 30'h0;
  assign io_covSum = Queue_15_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[6:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLError(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [3:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_corrupt,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  a_clock; // @[Decoupled.scala 361:21]
  wire  a_reset; // @[Decoupled.scala 361:21]
  wire  a_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  a_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] a_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] a_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] a_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire  a_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  a_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] a_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] a_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] a_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [29:0] a_io_covSum; // @[Decoupled.scala 361:21]
  wire  _a_last_T = a_io_deq_ready & a_io_deq_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _a_last_beats1_decode_T_1 = 27'hfff << a_io_deq_bits_size; // @[package.scala 234:77]
  wire [11:0] _a_last_beats1_decode_T_3 = ~_a_last_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] a_last_beats1_decode = _a_last_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  a_last_beats1_opdata = ~a_io_deq_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [8:0] a_last_beats1 = a_last_beats1_opdata ? a_last_beats1_decode : 9'h0; // @[Edges.scala 220:14]
  reg [8:0] a_last_counter; // @[Edges.scala 228:27]
  wire [8:0] a_last_counter1 = a_last_counter - 9'h1; // @[Edges.scala 229:28]
  wire  a_last_first = a_last_counter == 9'h0; // @[Edges.scala 230:25]
  wire  a_last = a_last_counter == 9'h1 | a_last_beats1 == 9'h0; // @[Edges.scala 231:37]
  wire  da_valid = a_io_deq_valid & a_last; // @[Error.scala 51:25]
  wire  _T = auto_in_d_ready & da_valid; // @[Decoupled.scala 50:35]
  wire [3:0] da_bits_size = a_io_deq_bits_size; // @[Error.scala 43:18 55:21]
  wire [26:0] _beats1_decode_T_1 = 27'hfff << da_bits_size; // @[package.scala 234:77]
  wire [11:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] beats1_decode = _beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire [2:0] _GEN_4 = 3'h2 == a_io_deq_bits_opcode ? 3'h1 : 3'h0; // @[Error.scala 53:{21,21}]
  wire [2:0] _GEN_5 = 3'h3 == a_io_deq_bits_opcode ? 3'h1 : _GEN_4; // @[Error.scala 53:{21,21}]
  wire [2:0] _GEN_6 = 3'h4 == a_io_deq_bits_opcode ? 3'h1 : _GEN_5; // @[Error.scala 53:{21,21}]
  wire [2:0] _GEN_7 = 3'h5 == a_io_deq_bits_opcode ? 3'h2 : _GEN_6; // @[Error.scala 53:{21,21}]
  wire [2:0] _GEN_8 = 3'h6 == a_io_deq_bits_opcode ? 3'h4 : _GEN_7; // @[Error.scala 53:{21,21}]
  wire [2:0] da_bits_opcode = 3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8; // @[Error.scala 53:{21,21}]
  wire  beats1_opdata = da_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [8:0] beats1 = beats1_opdata ? beats1_decode : 9'h0; // @[Edges.scala 220:14]
  reg [8:0] counter; // @[Edges.scala 228:27]
  wire [8:0] counter1 = counter - 9'h1; // @[Edges.scala 229:28]
  wire  da_first = counter == 9'h0; // @[Edges.scala 230:25]
  wire  da_last = counter == 9'h1 | beats1 == 9'h0; // @[Edges.scala 231:37]
  wire [29:0] TLError_covSum;
  wire [29:0] a_sum;
  Queue_15 a ( // @[Decoupled.scala 361:21]
    .clock(a_clock),
    .reset(a_reset),
    .io_enq_ready(a_io_enq_ready),
    .io_enq_valid(a_io_enq_valid),
    .io_enq_bits_opcode(a_io_enq_bits_opcode),
    .io_enq_bits_size(a_io_enq_bits_size),
    .io_enq_bits_source(a_io_enq_bits_source),
    .io_deq_ready(a_io_deq_ready),
    .io_deq_valid(a_io_deq_valid),
    .io_deq_bits_opcode(a_io_deq_bits_opcode),
    .io_deq_bits_size(a_io_deq_bits_size),
    .io_deq_bits_source(a_io_deq_bits_source),
    .io_covSum(a_io_covSum)
  );
  assign auto_in_a_ready = a_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_d_valid = a_io_deq_valid & a_last; // @[Error.scala 51:25]
  assign auto_in_d_bits_opcode = 3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8; // @[Error.scala 53:{21,21}]
  assign auto_in_d_bits_size = a_io_deq_bits_size; // @[Error.scala 43:18 55:21]
  assign auto_in_d_bits_source = a_io_deq_bits_source; // @[Error.scala 43:18 56:21]
  assign auto_in_d_bits_corrupt = da_bits_opcode[0]; // @[Edges.scala 105:36]
  assign a_clock = clock;
  assign a_reset = reset;
  assign a_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign a_io_deq_ready = auto_in_d_ready & da_last | ~a_last; // @[Error.scala 50:46]
  assign TLError_covSum = 30'h0;
  assign a_sum = TLError_covSum + a_io_covSum;
  assign io_covSum = a_sum;
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_last_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_a_last_T) begin
      if (a_last_first) begin
        if (a_last_beats1_opdata) begin
          a_last_counter <= a_last_beats1_decode;
        end else begin
          a_last_counter <= 9'h0;
        end
      end else begin
        a_last_counter <= a_last_counter1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_T) begin
      if (da_first) begin
        if (beats1_opdata) begin
          counter <= beats1_decode;
        end else begin
          counter <= 9'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Error.scala 49:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_last_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_16(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [3:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [3:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [6:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_16_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_16_covSum = 30'h0;
  assign io_covSum = Queue_16_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= value_1 + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[6:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_5(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [3:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [3:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum
);
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [29:0] bundleOut_0_a_q_io_covSum; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [6:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire [29:0] bundleIn_0_d_q_io_covSum; // @[Decoupled.scala 361:21]
  wire [29:0] TLBuffer_5_covSum;
  wire [29:0] bundleOut_0_a_q_sum;
  wire [29:0] bundleIn_0_d_q_sum;
  Queue_16 bundleOut_0_a_q ( // @[Decoupled.scala 361:21]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_covSum(bundleOut_0_a_q_io_covSum)
  );
  Queue_14 bundleIn_0_d_q ( // @[Decoupled.scala 361:21]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt),
    .io_covSum(bundleIn_0_d_q_io_covSum)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 Decoupled.scala 365:17]
  assign bundleOut_0_a_q_clock = clock;
  assign bundleOut_0_a_q_reset = reset;
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_clock = clock;
  assign bundleIn_0_d_q_reset = reset;
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_denied = 1'h1; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_data = 64'h0; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBuffer_5_covSum = 30'h0;
  assign bundleOut_0_a_q_sum = TLBuffer_5_covSum + bundleOut_0_a_q_io_covSum;
  assign bundleIn_0_d_q_sum = bundleOut_0_a_q_sum + bundleIn_0_d_q_io_covSum;
  assign io_covSum = bundleIn_0_d_q_sum;
endmodule
module ErrorDeviceWrapper(
  input         clock,
  input         reset,
  output        auto_buffer_in_a_ready,
  input         auto_buffer_in_a_valid,
  input  [2:0]  auto_buffer_in_a_bits_opcode,
  input  [3:0]  auto_buffer_in_a_bits_size,
  input  [6:0]  auto_buffer_in_a_bits_source,
  input         auto_buffer_in_d_ready,
  output        auto_buffer_in_d_valid,
  output [2:0]  auto_buffer_in_d_bits_opcode,
  output [3:0]  auto_buffer_in_d_bits_size,
  output [6:0]  auto_buffer_in_d_bits_source,
  output        auto_buffer_in_d_bits_denied,
  output [63:0] auto_buffer_in_d_bits_data,
  output        auto_buffer_in_d_bits_corrupt,
  output [29:0] io_covSum
);
  wire  error_clock; // @[CanHaveBuiltInDevices.scala 38:29]
  wire  error_reset; // @[CanHaveBuiltInDevices.scala 38:29]
  wire  error_auto_in_a_ready; // @[CanHaveBuiltInDevices.scala 38:29]
  wire  error_auto_in_a_valid; // @[CanHaveBuiltInDevices.scala 38:29]
  wire [2:0] error_auto_in_a_bits_opcode; // @[CanHaveBuiltInDevices.scala 38:29]
  wire [3:0] error_auto_in_a_bits_size; // @[CanHaveBuiltInDevices.scala 38:29]
  wire [6:0] error_auto_in_a_bits_source; // @[CanHaveBuiltInDevices.scala 38:29]
  wire  error_auto_in_d_ready; // @[CanHaveBuiltInDevices.scala 38:29]
  wire  error_auto_in_d_valid; // @[CanHaveBuiltInDevices.scala 38:29]
  wire [2:0] error_auto_in_d_bits_opcode; // @[CanHaveBuiltInDevices.scala 38:29]
  wire [3:0] error_auto_in_d_bits_size; // @[CanHaveBuiltInDevices.scala 38:29]
  wire [6:0] error_auto_in_d_bits_source; // @[CanHaveBuiltInDevices.scala 38:29]
  wire  error_auto_in_d_bits_corrupt; // @[CanHaveBuiltInDevices.scala 38:29]
  wire [29:0] error_io_covSum; // @[CanHaveBuiltInDevices.scala 38:29]
  wire  buffer_clock; // @[Buffer.scala 68:28]
  wire  buffer_reset; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire [29:0] buffer_io_covSum; // @[Buffer.scala 68:28]
  wire [29:0] ErrorDeviceWrapper_covSum;
  wire [29:0] error_sum;
  wire [29:0] buffer_sum;
  TLError error ( // @[CanHaveBuiltInDevices.scala 38:29]
    .clock(error_clock),
    .reset(error_reset),
    .auto_in_a_ready(error_auto_in_a_ready),
    .auto_in_a_valid(error_auto_in_a_valid),
    .auto_in_a_bits_opcode(error_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(error_auto_in_a_bits_size),
    .auto_in_a_bits_source(error_auto_in_a_bits_source),
    .auto_in_d_ready(error_auto_in_d_ready),
    .auto_in_d_valid(error_auto_in_d_valid),
    .auto_in_d_bits_opcode(error_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(error_auto_in_d_bits_size),
    .auto_in_d_bits_source(error_auto_in_d_bits_source),
    .auto_in_d_bits_corrupt(error_auto_in_d_bits_corrupt),
    .io_covSum(error_io_covSum)
  );
  TLBuffer_5 buffer ( // @[Buffer.scala 68:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt),
    .io_covSum(buffer_io_covSum)
  );
  assign auto_buffer_in_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 309:16]
  assign auto_buffer_in_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 309:16]
  assign auto_buffer_in_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign auto_buffer_in_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_buffer_in_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign auto_buffer_in_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 309:16]
  assign auto_buffer_in_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign auto_buffer_in_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign error_clock = clock;
  assign error_reset = reset;
  assign error_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign error_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign error_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign error_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign error_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_a_valid = auto_buffer_in_a_valid; // @[LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_opcode = auto_buffer_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_size = auto_buffer_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_source = auto_buffer_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign buffer_auto_in_d_ready = auto_buffer_in_d_ready; // @[LazyModule.scala 309:16]
  assign buffer_auto_out_a_ready = error_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_valid = error_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_opcode = error_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_size = error_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_source = error_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_corrupt = error_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign ErrorDeviceWrapper_covSum = 30'h0;
  assign error_sum = ErrorDeviceWrapper_covSum + error_io_covSum;
  assign buffer_sum = error_sum + buffer_io_covSum;
  assign io_covSum = buffer_sum;
endmodule
module Repeater_1(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [27:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [27:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [6:0] saved_source; // @[Repeater.scala 20:18]
  reg [27:0] saved_address; // @[Repeater.scala 20:18]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 19:21 28:{38,45}]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  reg  Repeater_1_covState; // @[Register tracking Repeater_1 state]
  reg  Repeater_1_covMap [0:1]; // @[Coverage map for Repeater_1]
  wire  Repeater_1_covMap_read_en; // @[Coverage map for Repeater_1]
  wire  Repeater_1_covMap_read_addr; // @[Coverage map for Repeater_1]
  wire  Repeater_1_covMap_read_data; // @[Coverage map for Repeater_1]
  wire  Repeater_1_covMap_write_data; // @[Coverage map for Repeater_1]
  wire  Repeater_1_covMap_write_addr; // @[Coverage map for Repeater_1]
  wire  Repeater_1_covMap_write_mask; // @[Coverage map for Repeater_1]
  wire  Repeater_1_covMap_write_en; // @[Coverage map for Repeater_1]
  reg [29:0] Repeater_1_covSum; // @[Sum of coverage map]
  wire  full_shl;
  wire  full_pad;
  assign io_full = full; // @[Repeater.scala 26:11]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21]
  assign Repeater_1_covMap_read_en = 1'h1;
  assign Repeater_1_covMap_read_addr = Repeater_1_covState;
  assign Repeater_1_covMap_read_data = Repeater_1_covMap[Repeater_1_covMap_read_addr]; // @[Coverage map for Repeater_1]
  assign Repeater_1_covMap_write_data = 1'h1;
  assign Repeater_1_covMap_write_addr = Repeater_1_covState;
  assign Repeater_1_covMap_write_mask = 1'h1;
  assign Repeater_1_covMap_write_en = ~metaReset;
  assign full_shl = full;
  assign full_pad = full_shl;
  assign io_covSum = Repeater_1_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin
      full <= 1'h0;
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62]
    end
    Repeater_1_covState <= full_pad;
    if (Repeater_1_covMap_write_en & Repeater_1_covMap_write_mask) begin
      Repeater_1_covMap[Repeater_1_covMap_write_addr] <= Repeater_1_covMap_write_data; // @[Coverage map for Repeater_1]
    end
    if (!(Repeater_1_covMap_read_data | metaReset)) begin
      Repeater_1_covSum <= Repeater_1_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Repeater_1_covMap[initvar] = 0; //_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_source = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  saved_address = _RAND_4[27:0];
  _RAND_5 = {1{`RANDOM}};
  saved_mask = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  Repeater_1_covState = 0; //_6[0:0];
  _RAND_8 = {1{`RANDOM}};
  Repeater_1_covSum = 0; //_8[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_1(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [27:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [1:0]  auto_out_a_bits_size,
  output [10:0] auto_out_a_bits_source,
  output [27:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_size,
  input  [10:0] auto_out_d_bits_source,
  input  [63:0] auto_out_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  repeater_clock; // @[Fragmenter.scala 262:30]
  wire  repeater_reset; // @[Fragmenter.scala 262:30]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_opcode; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30]
  wire [27:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_opcode; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30]
  wire [27:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30]
  wire [29:0] repeater_io_covSum; // @[Fragmenter.scala 262:30]
  wire  repeater_metaReset; // @[Fragmenter.scala 262:30]
  reg [2:0] acknum; // @[Fragmenter.scala 189:29]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24]
  reg  dToggle; // @[Fragmenter.scala 191:30]
  wire [2:0] dFragnum = auto_out_d_bits_source[2:0]; // @[Fragmenter.scala 192:41]
  wire  dFirst = acknum == 3'h0; // @[Fragmenter.scala 193:29]
  wire  dLast = dFragnum == 3'h0; // @[Fragmenter.scala 194:30]
  wire [3:0] dsizeOH = 4'h1 << auto_out_d_bits_size; // @[OneHot.scala 64:12]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[package.scala 234:46]
  wire  dHasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  _T_5 = ~reset; // @[Fragmenter.scala 202:16]
  wire  ack_decrement = dHasData | dsizeOH[3]; // @[Fragmenter.scala 204:32]
  wire [5:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[Fragmenter.scala 206:47]
  wire [5:0] _GEN_7 = {{3'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69]
  wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69]
  wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0}; // @[package.scala 232:35]
  wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h1; // @[package.scala 232:40]
  wire [6:0] _dFirst_size_T_4 = {1'h0,_dFirst_size_T_1}; // @[Cat.scala 31:58]
  wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4; // @[package.scala 232:53]
  wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5; // @[package.scala 232:51]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4]; // @[OneHot.scala 30:18]
  wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_7 = |dFirst_size_hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28]
  wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo; // @[OneHot.scala 32:28]
  wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_9 = |dFirst_size_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] dFirst_size = {_dFirst_size_T_7,_dFirst_size_T_9,_dFirst_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  drop = ~dHasData & ~dLast; // @[Fragmenter.scala 222:30]
  wire  bundleOut_0_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35]
  wire  _T_7 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_9 = {{2'd0}, ack_decrement}; // @[Fragmenter.scala 209:55]
  wire [2:0] _acknum_T_1 = acknum - _GEN_9; // @[Fragmenter.scala 209:55]
  wire [2:0] aFrag = repeater_io_deq_bits_size > 3'h3 ? 3'h3 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[package.scala 234:77]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[package.scala 234:46]
  wire  aHasData = ~repeater_io_deq_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] gennum; // @[Fragmenter.scala 291:29]
  wire  aFirst = gennum == 3'h0; // @[Fragmenter.scala 292:29]
  wire [2:0] _old_gennum1_T_2 = gennum - 3'h1; // @[Fragmenter.scala 293:79]
  wire [2:0] old_gennum1 = aFirst ? aOrigOH1[5:3] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30]
  wire [2:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28]
  wire [2:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26]
  reg  aToggle_r; // @[Reg.scala 16:16]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  aToggle = ~_GEN_5; // @[Fragmenter.scala 297:23]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 50:35]
  wire  _repeater_io_repeat_T = ~aHasData; // @[Fragmenter.scala 302:31]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 3'h0}; // @[Fragmenter.scala 304:65]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88]
  wire [5:0] _GEN_10 = {{3'd0}, aFragOH1}; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h7; // @[Fragmenter.scala 304:111]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51]
  wire [27:0] _GEN_11 = {{22'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49]
  wire [7:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,aToggle}; // @[Cat.scala 31:58]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17]
  wire [29:0] TLFragmenter_1_covSum;
  wire [29:0] repeater_sum;
  Repeater_1 repeater ( // @[Fragmenter.scala 262:30]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_opcode(repeater_io_enq_bits_opcode),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_opcode(repeater_io_deq_bits_opcode),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_covSum(repeater_io_covSum),
    .metaReset(repeater_metaReset)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 Fragmenter.scala 263:25]
  assign auto_in_d_valid = auto_out_d_valid & ~drop; // @[Fragmenter.scala 224:36]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32]
  assign auto_in_d_bits_source = auto_out_d_bits_source[10:4]; // @[Fragmenter.scala 226:47]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 Fragmenter.scala 306:25]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 31:58]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11; // @[Fragmenter.scala 304:49]
  assign auto_out_a_bits_mask = repeater_io_full ? 8'hff : auto_in_a_bits_mask; // @[Fragmenter.scala 313:31]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35]
  assign repeater_clock = clock;
  assign repeater_reset = reset;
  assign repeater_io_repeat = ~aHasData & new_gennum != 3'h0; // @[Fragmenter.scala 302:41]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign TLFragmenter_1_covSum = 30'h0;
  assign repeater_sum = TLFragmenter_1_covSum + repeater_io_covSum;
  assign io_covSum = repeater_sum;
  assign repeater_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29]
      acknum <= 3'h0; // @[Fragmenter.scala 189:29]
    end else if (_T_7) begin
      if (dFirst) begin
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29]
      if (dFirst) begin
        dOrig <= dFirst_size;
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30]
    end else if (_T_7) begin
      if (dFirst) begin
        dToggle <= auto_out_d_bits_source[3];
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29]
      gennum <= 3'h0; // @[Fragmenter.scala 291:29]
    end else if (_T_8) begin
      gennum <= new_gennum;
    end
    if (aFirst) begin // @[Reg.scala 17:18]
      aToggle_r <= dToggle; // @[Reg.scala 17:22]
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Fragmenter.scala 202:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~repeater_io_full | _repeater_io_repeat_T) & _T_5) begin
          $fatal; // @[Fragmenter.scala 309:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(~repeater_io_full | _repeater_io_repeat_T)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:309 assert (!repeater.io.full || !aHasData)\n"
            ); // @[Fragmenter.scala 309:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_9 | repeater_io_deq_bits_mask == 8'hff) & _T_5) begin
          $fatal; // @[Fragmenter.scala 312:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(_T_9 | repeater_io_deq_bits_mask == 8'hff)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLInterconnectCoupler_7(
  input         clock,
  input         reset,
  input         auto_fragmenter_out_a_ready,
  output        auto_fragmenter_out_a_valid,
  output [2:0]  auto_fragmenter_out_a_bits_opcode,
  output [1:0]  auto_fragmenter_out_a_bits_size,
  output [10:0] auto_fragmenter_out_a_bits_source,
  output [27:0] auto_fragmenter_out_a_bits_address,
  output [7:0]  auto_fragmenter_out_a_bits_mask,
  output [63:0] auto_fragmenter_out_a_bits_data,
  output        auto_fragmenter_out_d_ready,
  input         auto_fragmenter_out_d_valid,
  input  [2:0]  auto_fragmenter_out_d_bits_opcode,
  input  [1:0]  auto_fragmenter_out_d_bits_size,
  input  [10:0] auto_fragmenter_out_d_bits_source,
  input  [63:0] auto_fragmenter_out_d_bits_data,
  output        auto_tl_in_a_ready,
  input         auto_tl_in_a_valid,
  input  [2:0]  auto_tl_in_a_bits_opcode,
  input  [2:0]  auto_tl_in_a_bits_size,
  input  [6:0]  auto_tl_in_a_bits_source,
  input  [27:0] auto_tl_in_a_bits_address,
  input  [7:0]  auto_tl_in_a_bits_mask,
  input  [63:0] auto_tl_in_a_bits_data,
  input         auto_tl_in_d_ready,
  output        auto_tl_in_d_valid,
  output [2:0]  auto_tl_in_d_bits_opcode,
  output [2:0]  auto_tl_in_d_bits_size,
  output [6:0]  auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [27:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_in_a_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_out_a_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [27:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [7:0] fragmenter_auto_out_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_out_a_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_out_d_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34]
  wire [29:0] fragmenter_io_covSum; // @[Fragmenter.scala 333:34]
  wire  fragmenter_metaReset; // @[Fragmenter.scala 333:34]
  wire [29:0] TLInterconnectCoupler_7_covSum;
  wire [29:0] fragmenter_sum;
  TLFragmenter_1 fragmenter ( // @[Fragmenter.scala 333:34]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .io_covSum(fragmenter_io_covSum),
    .metaReset(fragmenter_metaReset)
  );
  assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_mask = fragmenter_auto_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_data = fragmenter_auto_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_opcode = fragmenter_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign fragmenter_clock = clock;
  assign fragmenter_reset = reset;
  assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_data = auto_tl_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_opcode = auto_fragmenter_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign TLInterconnectCoupler_7_covSum = 30'h0;
  assign fragmenter_sum = TLInterconnectCoupler_7_covSum + fragmenter_io_covSum;
  assign io_covSum = fragmenter_sum;
  assign fragmenter_metaReset = metaReset;
endmodule
module Repeater_2(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [25:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [25:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [6:0] saved_source; // @[Repeater.scala 20:18]
  reg [25:0] saved_address; // @[Repeater.scala 20:18]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 19:21 28:{38,45}]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  reg  Repeater_2_covState; // @[Register tracking Repeater_2 state]
  reg  Repeater_2_covMap [0:1]; // @[Coverage map for Repeater_2]
  wire  Repeater_2_covMap_read_en; // @[Coverage map for Repeater_2]
  wire  Repeater_2_covMap_read_addr; // @[Coverage map for Repeater_2]
  wire  Repeater_2_covMap_read_data; // @[Coverage map for Repeater_2]
  wire  Repeater_2_covMap_write_data; // @[Coverage map for Repeater_2]
  wire  Repeater_2_covMap_write_addr; // @[Coverage map for Repeater_2]
  wire  Repeater_2_covMap_write_mask; // @[Coverage map for Repeater_2]
  wire  Repeater_2_covMap_write_en; // @[Coverage map for Repeater_2]
  reg [29:0] Repeater_2_covSum; // @[Sum of coverage map]
  wire  full_shl;
  wire  full_pad;
  assign io_full = full; // @[Repeater.scala 26:11]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21]
  assign Repeater_2_covMap_read_en = 1'h1;
  assign Repeater_2_covMap_read_addr = Repeater_2_covState;
  assign Repeater_2_covMap_read_data = Repeater_2_covMap[Repeater_2_covMap_read_addr]; // @[Coverage map for Repeater_2]
  assign Repeater_2_covMap_write_data = 1'h1;
  assign Repeater_2_covMap_write_addr = Repeater_2_covState;
  assign Repeater_2_covMap_write_mask = 1'h1;
  assign Repeater_2_covMap_write_en = ~metaReset;
  assign full_shl = full;
  assign full_pad = full_shl;
  assign io_covSum = Repeater_2_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin
      full <= 1'h0;
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62]
    end
    Repeater_2_covState <= full_pad;
    if (Repeater_2_covMap_write_en & Repeater_2_covMap_write_mask) begin
      Repeater_2_covMap[Repeater_2_covMap_write_addr] <= Repeater_2_covMap_write_data; // @[Coverage map for Repeater_2]
    end
    if (!(Repeater_2_covMap_read_data | metaReset)) begin
      Repeater_2_covSum <= Repeater_2_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Repeater_2_covMap[initvar] = 0; //_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_source = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  saved_address = _RAND_4[25:0];
  _RAND_5 = {1{`RANDOM}};
  saved_mask = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  Repeater_2_covState = 0; //_6[0:0];
  _RAND_8 = {1{`RANDOM}};
  Repeater_2_covSum = 0; //_8[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_2(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [25:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [1:0]  auto_out_a_bits_size,
  output [10:0] auto_out_a_bits_source,
  output [25:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_size,
  input  [10:0] auto_out_d_bits_source,
  input  [63:0] auto_out_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  repeater_clock; // @[Fragmenter.scala 262:30]
  wire  repeater_reset; // @[Fragmenter.scala 262:30]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_opcode; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30]
  wire [25:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_opcode; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30]
  wire [25:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30]
  wire [29:0] repeater_io_covSum; // @[Fragmenter.scala 262:30]
  wire  repeater_metaReset; // @[Fragmenter.scala 262:30]
  reg [2:0] acknum; // @[Fragmenter.scala 189:29]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24]
  reg  dToggle; // @[Fragmenter.scala 191:30]
  wire [2:0] dFragnum = auto_out_d_bits_source[2:0]; // @[Fragmenter.scala 192:41]
  wire  dFirst = acknum == 3'h0; // @[Fragmenter.scala 193:29]
  wire  dLast = dFragnum == 3'h0; // @[Fragmenter.scala 194:30]
  wire [3:0] dsizeOH = 4'h1 << auto_out_d_bits_size; // @[OneHot.scala 64:12]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[package.scala 234:46]
  wire  dHasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  _T_5 = ~reset; // @[Fragmenter.scala 202:16]
  wire  ack_decrement = dHasData | dsizeOH[3]; // @[Fragmenter.scala 204:32]
  wire [5:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[Fragmenter.scala 206:47]
  wire [5:0] _GEN_7 = {{3'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69]
  wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69]
  wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0}; // @[package.scala 232:35]
  wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h1; // @[package.scala 232:40]
  wire [6:0] _dFirst_size_T_4 = {1'h0,_dFirst_size_T_1}; // @[Cat.scala 31:58]
  wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4; // @[package.scala 232:53]
  wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5; // @[package.scala 232:51]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4]; // @[OneHot.scala 30:18]
  wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_7 = |dFirst_size_hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28]
  wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo; // @[OneHot.scala 32:28]
  wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_9 = |dFirst_size_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] dFirst_size = {_dFirst_size_T_7,_dFirst_size_T_9,_dFirst_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  drop = ~dHasData & ~dLast; // @[Fragmenter.scala 222:30]
  wire  bundleOut_0_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35]
  wire  _T_7 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_9 = {{2'd0}, ack_decrement}; // @[Fragmenter.scala 209:55]
  wire [2:0] _acknum_T_1 = acknum - _GEN_9; // @[Fragmenter.scala 209:55]
  wire [2:0] aFrag = repeater_io_deq_bits_size > 3'h3 ? 3'h3 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[package.scala 234:77]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[package.scala 234:46]
  wire  aHasData = ~repeater_io_deq_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] gennum; // @[Fragmenter.scala 291:29]
  wire  aFirst = gennum == 3'h0; // @[Fragmenter.scala 292:29]
  wire [2:0] _old_gennum1_T_2 = gennum - 3'h1; // @[Fragmenter.scala 293:79]
  wire [2:0] old_gennum1 = aFirst ? aOrigOH1[5:3] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30]
  wire [2:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28]
  wire [2:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26]
  reg  aToggle_r; // @[Reg.scala 16:16]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  aToggle = ~_GEN_5; // @[Fragmenter.scala 297:23]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 50:35]
  wire  _repeater_io_repeat_T = ~aHasData; // @[Fragmenter.scala 302:31]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 3'h0}; // @[Fragmenter.scala 304:65]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88]
  wire [5:0] _GEN_10 = {{3'd0}, aFragOH1}; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h7; // @[Fragmenter.scala 304:111]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51]
  wire [25:0] _GEN_11 = {{20'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49]
  wire [7:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,aToggle}; // @[Cat.scala 31:58]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17]
  wire [29:0] TLFragmenter_2_covSum;
  wire [29:0] repeater_sum;
  Repeater_2 repeater ( // @[Fragmenter.scala 262:30]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_opcode(repeater_io_enq_bits_opcode),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_opcode(repeater_io_deq_bits_opcode),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_covSum(repeater_io_covSum),
    .metaReset(repeater_metaReset)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 Fragmenter.scala 263:25]
  assign auto_in_d_valid = auto_out_d_valid & ~drop; // @[Fragmenter.scala 224:36]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32]
  assign auto_in_d_bits_source = auto_out_d_bits_source[10:4]; // @[Fragmenter.scala 226:47]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 Fragmenter.scala 306:25]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 31:58]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11; // @[Fragmenter.scala 304:49]
  assign auto_out_a_bits_mask = repeater_io_full ? 8'hff : auto_in_a_bits_mask; // @[Fragmenter.scala 313:31]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35]
  assign repeater_clock = clock;
  assign repeater_reset = reset;
  assign repeater_io_repeat = ~aHasData & new_gennum != 3'h0; // @[Fragmenter.scala 302:41]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign TLFragmenter_2_covSum = 30'h0;
  assign repeater_sum = TLFragmenter_2_covSum + repeater_io_covSum;
  assign io_covSum = repeater_sum;
  assign repeater_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29]
      acknum <= 3'h0; // @[Fragmenter.scala 189:29]
    end else if (_T_7) begin
      if (dFirst) begin
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29]
      if (dFirst) begin
        dOrig <= dFirst_size;
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30]
    end else if (_T_7) begin
      if (dFirst) begin
        dToggle <= auto_out_d_bits_source[3];
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29]
      gennum <= 3'h0; // @[Fragmenter.scala 291:29]
    end else if (_T_8) begin
      gennum <= new_gennum;
    end
    if (aFirst) begin // @[Reg.scala 17:18]
      aToggle_r <= dToggle; // @[Reg.scala 17:22]
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Fragmenter.scala 202:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~repeater_io_full | _repeater_io_repeat_T) & _T_5) begin
          $fatal; // @[Fragmenter.scala 309:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(~repeater_io_full | _repeater_io_repeat_T)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:309 assert (!repeater.io.full || !aHasData)\n"
            ); // @[Fragmenter.scala 309:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_9 | repeater_io_deq_bits_mask == 8'hff) & _T_5) begin
          $fatal; // @[Fragmenter.scala 312:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(_T_9 | repeater_io_deq_bits_mask == 8'hff)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLInterconnectCoupler_8(
  input         clock,
  input         reset,
  input         auto_fragmenter_out_a_ready,
  output        auto_fragmenter_out_a_valid,
  output [2:0]  auto_fragmenter_out_a_bits_opcode,
  output [1:0]  auto_fragmenter_out_a_bits_size,
  output [10:0] auto_fragmenter_out_a_bits_source,
  output [25:0] auto_fragmenter_out_a_bits_address,
  output [7:0]  auto_fragmenter_out_a_bits_mask,
  output [63:0] auto_fragmenter_out_a_bits_data,
  output        auto_fragmenter_out_d_ready,
  input         auto_fragmenter_out_d_valid,
  input  [2:0]  auto_fragmenter_out_d_bits_opcode,
  input  [1:0]  auto_fragmenter_out_d_bits_size,
  input  [10:0] auto_fragmenter_out_d_bits_source,
  input  [63:0] auto_fragmenter_out_d_bits_data,
  output        auto_tl_in_a_ready,
  input         auto_tl_in_a_valid,
  input  [2:0]  auto_tl_in_a_bits_opcode,
  input  [2:0]  auto_tl_in_a_bits_size,
  input  [6:0]  auto_tl_in_a_bits_source,
  input  [25:0] auto_tl_in_a_bits_address,
  input  [7:0]  auto_tl_in_a_bits_mask,
  input  [63:0] auto_tl_in_a_bits_data,
  input         auto_tl_in_d_ready,
  output        auto_tl_in_d_valid,
  output [2:0]  auto_tl_in_d_bits_opcode,
  output [2:0]  auto_tl_in_d_bits_size,
  output [6:0]  auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [25:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_in_a_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_out_a_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [25:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [7:0] fragmenter_auto_out_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_out_a_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_out_d_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34]
  wire [29:0] fragmenter_io_covSum; // @[Fragmenter.scala 333:34]
  wire  fragmenter_metaReset; // @[Fragmenter.scala 333:34]
  wire [29:0] TLInterconnectCoupler_8_covSum;
  wire [29:0] fragmenter_sum;
  TLFragmenter_2 fragmenter ( // @[Fragmenter.scala 333:34]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .io_covSum(fragmenter_io_covSum),
    .metaReset(fragmenter_metaReset)
  );
  assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_mask = fragmenter_auto_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_data = fragmenter_auto_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_opcode = fragmenter_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign fragmenter_clock = clock;
  assign fragmenter_reset = reset;
  assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_data = auto_tl_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_opcode = auto_fragmenter_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign TLInterconnectCoupler_8_covSum = 30'h0;
  assign fragmenter_sum = TLInterconnectCoupler_8_covSum + fragmenter_io_covSum;
  assign io_covSum = fragmenter_sum;
  assign fragmenter_metaReset = metaReset;
endmodule
module Repeater_3(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [16:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [16:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [6:0] saved_source; // @[Repeater.scala 20:18]
  reg [16:0] saved_address; // @[Repeater.scala 20:18]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 19:21 28:{38,45}]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  reg  Repeater_3_covState; // @[Register tracking Repeater_3 state]
  reg  Repeater_3_covMap [0:1]; // @[Coverage map for Repeater_3]
  wire  Repeater_3_covMap_read_en; // @[Coverage map for Repeater_3]
  wire  Repeater_3_covMap_read_addr; // @[Coverage map for Repeater_3]
  wire  Repeater_3_covMap_read_data; // @[Coverage map for Repeater_3]
  wire  Repeater_3_covMap_write_data; // @[Coverage map for Repeater_3]
  wire  Repeater_3_covMap_write_addr; // @[Coverage map for Repeater_3]
  wire  Repeater_3_covMap_write_mask; // @[Coverage map for Repeater_3]
  wire  Repeater_3_covMap_write_en; // @[Coverage map for Repeater_3]
  reg [29:0] Repeater_3_covSum; // @[Sum of coverage map]
  wire  full_shl;
  wire  full_pad;
  assign io_full = full; // @[Repeater.scala 26:11]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21]
  assign Repeater_3_covMap_read_en = 1'h1;
  assign Repeater_3_covMap_read_addr = Repeater_3_covState;
  assign Repeater_3_covMap_read_data = Repeater_3_covMap[Repeater_3_covMap_read_addr]; // @[Coverage map for Repeater_3]
  assign Repeater_3_covMap_write_data = 1'h1;
  assign Repeater_3_covMap_write_addr = Repeater_3_covState;
  assign Repeater_3_covMap_write_mask = 1'h1;
  assign Repeater_3_covMap_write_en = ~metaReset;
  assign full_shl = full;
  assign full_pad = full_shl;
  assign io_covSum = Repeater_3_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin
      full <= 1'h0;
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62]
    end
    Repeater_3_covState <= full_pad;
    if (Repeater_3_covMap_write_en & Repeater_3_covMap_write_mask) begin
      Repeater_3_covMap[Repeater_3_covMap_write_addr] <= Repeater_3_covMap_write_data; // @[Coverage map for Repeater_3]
    end
    if (!(Repeater_3_covMap_read_data | metaReset)) begin
      Repeater_3_covSum <= Repeater_3_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Repeater_3_covMap[initvar] = 0; //_6[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_size = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_source = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  saved_address = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  saved_mask = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  Repeater_3_covState = 0; //_5[0:0];
  _RAND_7 = {1{`RANDOM}};
  Repeater_3_covSum = 0; //_7[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_3(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [16:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [1:0]  auto_out_a_bits_size,
  output [10:0] auto_out_a_bits_source,
  output [16:0] auto_out_a_bits_address,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [1:0]  auto_out_d_bits_size,
  input  [10:0] auto_out_d_bits_source,
  input  [63:0] auto_out_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  repeater_clock; // @[Fragmenter.scala 262:30]
  wire  repeater_reset; // @[Fragmenter.scala 262:30]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30]
  wire [16:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30]
  wire [16:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30]
  wire [29:0] repeater_io_covSum; // @[Fragmenter.scala 262:30]
  wire  repeater_metaReset; // @[Fragmenter.scala 262:30]
  reg [2:0] acknum; // @[Fragmenter.scala 189:29]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24]
  reg  dToggle; // @[Fragmenter.scala 191:30]
  wire [2:0] dFragnum = auto_out_d_bits_source[2:0]; // @[Fragmenter.scala 192:41]
  wire  dFirst = acknum == 3'h0; // @[Fragmenter.scala 193:29]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[package.scala 234:46]
  wire  _T_5 = ~reset; // @[Fragmenter.scala 202:16]
  wire [5:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[Fragmenter.scala 206:47]
  wire [5:0] _GEN_7 = {{3'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69]
  wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69]
  wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0}; // @[package.scala 232:35]
  wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h1; // @[package.scala 232:40]
  wire [6:0] _dFirst_size_T_4 = {1'h0,_dFirst_size_T_1}; // @[Cat.scala 31:58]
  wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4; // @[package.scala 232:53]
  wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5; // @[package.scala 232:51]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4]; // @[OneHot.scala 30:18]
  wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_7 = |dFirst_size_hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28]
  wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo; // @[OneHot.scala 32:28]
  wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_9 = |dFirst_size_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] dFirst_size = {_dFirst_size_T_7,_dFirst_size_T_9,_dFirst_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  _T_7 = auto_in_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _acknum_T_1 = acknum - 3'h1; // @[Fragmenter.scala 209:55]
  wire [2:0] aFrag = repeater_io_deq_bits_size > 3'h3 ? 3'h3 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[package.scala 234:77]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[package.scala 234:46]
  reg [2:0] gennum; // @[Fragmenter.scala 291:29]
  wire  aFirst = gennum == 3'h0; // @[Fragmenter.scala 292:29]
  wire [2:0] _old_gennum1_T_2 = gennum - 3'h1; // @[Fragmenter.scala 293:79]
  wire [2:0] old_gennum1 = aFirst ? aOrigOH1[5:3] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30]
  wire [2:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28]
  wire [2:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26]
  reg  aToggle_r; // @[Reg.scala 16:16]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  aToggle = ~_GEN_5; // @[Fragmenter.scala 297:23]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 3'h0}; // @[Fragmenter.scala 304:65]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88]
  wire [5:0] _GEN_9 = {{3'd0}, aFragOH1}; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_9; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h7; // @[Fragmenter.scala 304:111]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51]
  wire [16:0] _GEN_10 = {{11'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49]
  wire [7:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,aToggle}; // @[Cat.scala 31:58]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17]
  wire [29:0] TLFragmenter_3_covSum;
  wire [29:0] repeater_sum;
  Repeater_3 repeater ( // @[Fragmenter.scala 262:30]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_covSum(repeater_io_covSum),
    .metaReset(repeater_metaReset)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 Fragmenter.scala 263:25]
  assign auto_in_d_valid = auto_out_d_valid; // @[Fragmenter.scala 224:36]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32]
  assign auto_in_d_bits_source = auto_out_d_bits_source[10:4]; // @[Fragmenter.scala 226:47]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 Fragmenter.scala 306:25]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 31:58]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_10; // @[Fragmenter.scala 304:49]
  assign auto_out_d_ready = auto_in_d_ready; // @[Fragmenter.scala 223:35]
  assign repeater_clock = clock;
  assign repeater_reset = reset;
  assign repeater_io_repeat = new_gennum != 3'h0; // @[Fragmenter.scala 302:53]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign TLFragmenter_3_covSum = 30'h0;
  assign repeater_sum = TLFragmenter_3_covSum + repeater_io_covSum;
  assign io_covSum = repeater_sum;
  assign repeater_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29]
      acknum <= 3'h0; // @[Fragmenter.scala 189:29]
    end else if (_T_7) begin
      if (dFirst) begin
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29]
      if (dFirst) begin
        dOrig <= dFirst_size;
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30]
    end else if (_T_7) begin
      if (dFirst) begin
        dToggle <= auto_out_d_bits_source[3];
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29]
      gennum <= 3'h0; // @[Fragmenter.scala 291:29]
    end else if (_T_8) begin
      gennum <= new_gennum;
    end
    if (aFirst) begin // @[Reg.scala 17:18]
      aToggle_r <= dToggle; // @[Reg.scala 17:22]
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Fragmenter.scala 202:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & _T_5) begin
          $fatal; // @[Fragmenter.scala 309:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_9 | repeater_io_deq_bits_mask == 8'hff) & _T_5) begin
          $fatal; // @[Fragmenter.scala 312:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(_T_9 | repeater_io_deq_bits_mask == 8'hff)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLInterconnectCoupler_10(
  input         clock,
  input         reset,
  input         auto_fragmenter_out_a_ready,
  output        auto_fragmenter_out_a_valid,
  output [1:0]  auto_fragmenter_out_a_bits_size,
  output [10:0] auto_fragmenter_out_a_bits_source,
  output [16:0] auto_fragmenter_out_a_bits_address,
  output        auto_fragmenter_out_d_ready,
  input         auto_fragmenter_out_d_valid,
  input  [1:0]  auto_fragmenter_out_d_bits_size,
  input  [10:0] auto_fragmenter_out_d_bits_source,
  input  [63:0] auto_fragmenter_out_d_bits_data,
  output        auto_tl_in_a_ready,
  input         auto_tl_in_a_valid,
  input  [2:0]  auto_tl_in_a_bits_size,
  input  [6:0]  auto_tl_in_a_bits_source,
  input  [16:0] auto_tl_in_a_bits_address,
  input  [7:0]  auto_tl_in_a_bits_mask,
  input         auto_tl_in_d_ready,
  output        auto_tl_in_d_valid,
  output [2:0]  auto_tl_in_d_bits_size,
  output [6:0]  auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [16:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [16:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34]
  wire [29:0] fragmenter_io_covSum; // @[Fragmenter.scala 333:34]
  wire  fragmenter_metaReset; // @[Fragmenter.scala 333:34]
  wire [29:0] TLInterconnectCoupler_10_covSum;
  wire [29:0] fragmenter_sum;
  TLFragmenter_3 fragmenter ( // @[Fragmenter.scala 333:34]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .io_covSum(fragmenter_io_covSum),
    .metaReset(fragmenter_metaReset)
  );
  assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign fragmenter_clock = clock;
  assign fragmenter_reset = reset;
  assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign TLInterconnectCoupler_10_covSum = 30'h0;
  assign fragmenter_sum = TLInterconnectCoupler_10_covSum + fragmenter_io_covSum;
  assign io_covSum = fragmenter_sum;
  assign fragmenter_metaReset = metaReset;
endmodule
module Repeater_4(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [17:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [17:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [6:0] saved_source; // @[Repeater.scala 20:18]
  reg [17:0] saved_address; // @[Repeater.scala 20:18]
  reg [3:0] saved_mask; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 19:21 28:{38,45}]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  reg  Repeater_4_covState; // @[Register tracking Repeater_4 state]
  reg  Repeater_4_covMap [0:1]; // @[Coverage map for Repeater_4]
  wire  Repeater_4_covMap_read_en; // @[Coverage map for Repeater_4]
  wire  Repeater_4_covMap_read_addr; // @[Coverage map for Repeater_4]
  wire  Repeater_4_covMap_read_data; // @[Coverage map for Repeater_4]
  wire  Repeater_4_covMap_write_data; // @[Coverage map for Repeater_4]
  wire  Repeater_4_covMap_write_addr; // @[Coverage map for Repeater_4]
  wire  Repeater_4_covMap_write_mask; // @[Coverage map for Repeater_4]
  wire  Repeater_4_covMap_write_en; // @[Coverage map for Repeater_4]
  reg [29:0] Repeater_4_covSum; // @[Sum of coverage map]
  wire  full_shl;
  wire  full_pad;
  assign io_full = full; // @[Repeater.scala 26:11]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21]
  assign Repeater_4_covMap_read_en = 1'h1;
  assign Repeater_4_covMap_read_addr = Repeater_4_covState;
  assign Repeater_4_covMap_read_data = Repeater_4_covMap[Repeater_4_covMap_read_addr]; // @[Coverage map for Repeater_4]
  assign Repeater_4_covMap_write_data = 1'h1;
  assign Repeater_4_covMap_write_addr = Repeater_4_covState;
  assign Repeater_4_covMap_write_mask = 1'h1;
  assign Repeater_4_covMap_write_en = ~metaReset;
  assign full_shl = full;
  assign full_pad = full_shl;
  assign io_covSum = Repeater_4_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin
      full <= 1'h0;
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62]
    end
    Repeater_4_covState <= full_pad;
    if (Repeater_4_covMap_write_en & Repeater_4_covMap_write_mask) begin
      Repeater_4_covMap[Repeater_4_covMap_write_addr] <= Repeater_4_covMap_write_data; // @[Coverage map for Repeater_4]
    end
    if (!(Repeater_4_covMap_read_data | metaReset)) begin
      Repeater_4_covSum <= Repeater_4_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Repeater_4_covMap[initvar] = 0; //_6[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_size = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_source = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  saved_address = _RAND_3[17:0];
  _RAND_4 = {1{`RANDOM}};
  saved_mask = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  Repeater_4_covState = 0; //_5[0:0];
  _RAND_7 = {1{`RANDOM}};
  Repeater_4_covSum = 0; //_7[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_4(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [17:0] auto_in_a_bits_address,
  input  [3:0]  auto_in_a_bits_mask,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output [31:0] auto_in_d_bits_data,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [1:0]  auto_out_a_bits_size,
  output [11:0] auto_out_a_bits_source,
  output [17:0] auto_out_a_bits_address,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [1:0]  auto_out_d_bits_size,
  input  [11:0] auto_out_d_bits_source,
  input  [31:0] auto_out_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  repeater_clock; // @[Fragmenter.scala 262:30]
  wire  repeater_reset; // @[Fragmenter.scala 262:30]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30]
  wire [17:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30]
  wire [3:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30]
  wire [17:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30]
  wire [3:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30]
  wire [29:0] repeater_io_covSum; // @[Fragmenter.scala 262:30]
  wire  repeater_metaReset; // @[Fragmenter.scala 262:30]
  reg [3:0] acknum; // @[Fragmenter.scala 189:29]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24]
  reg  dToggle; // @[Fragmenter.scala 191:30]
  wire [3:0] dFragnum = auto_out_d_bits_source[3:0]; // @[Fragmenter.scala 192:41]
  wire  dFirst = acknum == 4'h0; // @[Fragmenter.scala 193:29]
  wire [4:0] _dsizeOH1_T_1 = 5'h3 << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0]; // @[package.scala 234:46]
  wire  _T_5 = ~reset; // @[Fragmenter.scala 202:16]
  wire [5:0] _dFirst_size_T = {dFragnum, 2'h0}; // @[Fragmenter.scala 206:47]
  wire [5:0] _GEN_7 = {{4'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69]
  wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69]
  wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0}; // @[package.scala 232:35]
  wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h1; // @[package.scala 232:40]
  wire [6:0] _dFirst_size_T_4 = {1'h0,_dFirst_size_T_1}; // @[Cat.scala 31:58]
  wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4; // @[package.scala 232:53]
  wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5; // @[package.scala 232:51]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4]; // @[OneHot.scala 30:18]
  wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_7 = |dFirst_size_hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28]
  wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo; // @[OneHot.scala 32:28]
  wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_9 = |dFirst_size_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] dFirst_size = {_dFirst_size_T_7,_dFirst_size_T_9,_dFirst_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  _T_7 = auto_in_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _acknum_T_1 = acknum - 4'h1; // @[Fragmenter.scala 209:55]
  wire [2:0] aFrag = repeater_io_deq_bits_size > 3'h2 ? 3'h2 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46]
  wire [8:0] _aFragOH1_T_1 = 9'h3 << aFrag; // @[package.scala 234:77]
  wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0]; // @[package.scala 234:46]
  reg [3:0] gennum; // @[Fragmenter.scala 291:29]
  wire  aFirst = gennum == 4'h0; // @[Fragmenter.scala 292:29]
  wire [3:0] _old_gennum1_T_2 = gennum - 4'h1; // @[Fragmenter.scala 293:79]
  wire [3:0] old_gennum1 = aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30]
  wire [3:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28]
  wire [3:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26]
  reg  aToggle_r; // @[Reg.scala 16:16]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  aToggle = ~_GEN_5; // @[Fragmenter.scala 297:23]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0}; // @[Fragmenter.scala 304:65]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88]
  wire [5:0] _GEN_9 = {{4'd0}, aFragOH1}; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_9; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h3; // @[Fragmenter.scala 304:111]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51]
  wire [17:0] _GEN_10 = {{12'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49]
  wire [7:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,aToggle}; // @[Cat.scala 31:58]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17]
  wire [29:0] TLFragmenter_4_covSum;
  wire [29:0] repeater_sum;
  Repeater_4 repeater ( // @[Fragmenter.scala 262:30]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_covSum(repeater_io_covSum),
    .metaReset(repeater_metaReset)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 Fragmenter.scala 263:25]
  assign auto_in_d_valid = auto_out_d_valid; // @[Fragmenter.scala 224:36]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32]
  assign auto_in_d_bits_source = auto_out_d_bits_source[11:5]; // @[Fragmenter.scala 226:47]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 Fragmenter.scala 306:25]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 31:58]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_10; // @[Fragmenter.scala 304:49]
  assign auto_out_d_ready = auto_in_d_ready; // @[Fragmenter.scala 223:35]
  assign repeater_clock = clock;
  assign repeater_reset = reset;
  assign repeater_io_repeat = new_gennum != 4'h0; // @[Fragmenter.scala 302:53]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign TLFragmenter_4_covSum = 30'h0;
  assign repeater_sum = TLFragmenter_4_covSum + repeater_io_covSum;
  assign io_covSum = repeater_sum;
  assign repeater_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29]
      acknum <= 4'h0; // @[Fragmenter.scala 189:29]
    end else if (_T_7) begin
      if (dFirst) begin
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29]
      if (dFirst) begin
        dOrig <= dFirst_size;
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30]
    end else if (_T_7) begin
      if (dFirst) begin
        dToggle <= auto_out_d_bits_source[4];
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29]
      gennum <= 4'h0; // @[Fragmenter.scala 291:29]
    end else if (_T_8) begin
      gennum <= new_gennum;
    end
    if (aFirst) begin // @[Reg.scala 17:18]
      aToggle_r <= dToggle; // @[Reg.scala 17:22]
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Fragmenter.scala 202:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & _T_5) begin
          $fatal; // @[Fragmenter.scala 309:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_9 | repeater_io_deq_bits_mask == 4'hf) & _T_5) begin
          $fatal; // @[Fragmenter.scala 312:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(_T_9 | repeater_io_deq_bits_mask == 4'hf)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_5(
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [17:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [17:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [29:0] io_covSum
);
  wire [29:0] Repeater_5_covSum;
  assign io_enq_ready = io_deq_ready; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid; // @[Repeater.scala 23:32]
  assign io_deq_bits_size = io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = io_enq_bits_address; // @[Repeater.scala 25:21]
  assign io_deq_bits_mask = io_enq_bits_mask; // @[Repeater.scala 25:21]
  assign Repeater_5_covSum = 30'h0;
  assign io_covSum = Repeater_5_covSum;
endmodule
module TLWidthWidget_6(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [17:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_size,
  output [6:0]  auto_out_a_bits_source,
  output [17:0] auto_out_a_bits_address,
  output [3:0]  auto_out_a_bits_mask,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_size,
  input  [6:0]  auto_out_d_bits_source,
  input  [31:0] auto_out_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  repeated_repeater_io_enq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_size; // @[Repeater.scala 35:26]
  wire [6:0] repeated_repeater_io_enq_bits_source; // @[Repeater.scala 35:26]
  wire [17:0] repeated_repeater_io_enq_bits_address; // @[Repeater.scala 35:26]
  wire [7:0] repeated_repeater_io_enq_bits_mask; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_size; // @[Repeater.scala 35:26]
  wire [6:0] repeated_repeater_io_deq_bits_source; // @[Repeater.scala 35:26]
  wire [17:0] repeated_repeater_io_deq_bits_address; // @[Repeater.scala 35:26]
  wire [7:0] repeated_repeater_io_deq_bits_mask; // @[Repeater.scala 35:26]
  wire [29:0] repeated_repeater_io_covSum; // @[Repeater.scala 35:26]
  wire [17:0] cated_bits_address = repeated_repeater_io_deq_bits_address; // @[WidthWidget.scala 155:25 156:15]
  wire  repeat_sel = cated_bits_address[2]; // @[WidthWidget.scala 110:39]
  wire [7:0] cated_bits_mask = repeated_repeater_io_deq_bits_mask; // @[WidthWidget.scala 155:25 156:15]
  wire [3:0] repeat_bundleOut_0_a_bits_mask_mux_0 = cated_bits_mask[3:0]; // @[WidthWidget.scala 122:55]
  wire [3:0] repeat_bundleOut_0_a_bits_mask_mux_1 = cated_bits_mask[7:4]; // @[WidthWidget.scala 122:55]
  wire [9:0] _limit_T_1 = 10'h7 << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [2:0] _limit_T_3 = ~_limit_T_1[2:0]; // @[package.scala 234:46]
  wire  limit = _limit_T_3[2]; // @[WidthWidget.scala 32:47]
  reg  count; // @[WidthWidget.scala 34:27]
  wire  last = count == limit; // @[WidthWidget.scala 36:26]
  wire  enable_0 = ~(|(count & limit)); // @[WidthWidget.scala 37:47]
  wire  _bundleOut_0_d_ready_T = ~last; // @[WidthWidget.scala 70:32]
  wire  bundleOut_0_d_ready = auto_in_d_ready | ~last; // @[WidthWidget.scala 70:29]
  wire  _T = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  reg  bundleIn_0_d_bits_data_rdata_written_once; // @[WidthWidget.scala 56:41]
  wire  bundleIn_0_d_bits_data_masked_enable_0 = enable_0 | ~bundleIn_0_d_bits_data_rdata_written_once; // @[WidthWidget.scala 57:42]
  reg [31:0] bundleIn_0_d_bits_data_rdata_0; // @[WidthWidget.scala 60:24]
  wire [31:0] bundleIn_0_d_bits_data_mdata_0 = bundleIn_0_d_bits_data_masked_enable_0 ? auto_out_d_bits_data :
    bundleIn_0_d_bits_data_rdata_0; // @[WidthWidget.scala 62:88]
  wire  _GEN_8 = _T & _bundleOut_0_d_ready_T | bundleIn_0_d_bits_data_rdata_written_once; // @[WidthWidget.scala 63:35 64:30 56:41]
  reg [1:0] TLWidthWidget_6_covState; // @[Register tracking TLWidthWidget_6 state]
  reg  TLWidthWidget_6_covMap [0:3]; // @[Coverage map for TLWidthWidget_6]
  wire  TLWidthWidget_6_covMap_read_en; // @[Coverage map for TLWidthWidget_6]
  wire [1:0] TLWidthWidget_6_covMap_read_addr; // @[Coverage map for TLWidthWidget_6]
  wire  TLWidthWidget_6_covMap_read_data; // @[Coverage map for TLWidthWidget_6]
  wire  TLWidthWidget_6_covMap_write_data; // @[Coverage map for TLWidthWidget_6]
  wire [1:0] TLWidthWidget_6_covMap_write_addr; // @[Coverage map for TLWidthWidget_6]
  wire  TLWidthWidget_6_covMap_write_mask; // @[Coverage map for TLWidthWidget_6]
  wire  TLWidthWidget_6_covMap_write_en; // @[Coverage map for TLWidthWidget_6]
  reg [29:0] TLWidthWidget_6_covSum; // @[Sum of coverage map]
  wire  bundleIn_0_d_bits_data_rdata_written_once_shl;
  wire [1:0] bundleIn_0_d_bits_data_rdata_written_once_pad;
  wire [1:0] count_shl;
  wire [1:0] count_pad;
  wire [1:0] TLWidthWidget_6_xor0;
  wire [29:0] repeated_repeater_sum;
  Repeater_5 repeated_repeater ( // @[Repeater.scala 35:26]
    .io_enq_ready(repeated_repeater_io_enq_ready),
    .io_enq_valid(repeated_repeater_io_enq_valid),
    .io_enq_bits_size(repeated_repeater_io_enq_bits_size),
    .io_enq_bits_source(repeated_repeater_io_enq_bits_source),
    .io_enq_bits_address(repeated_repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeated_repeater_io_enq_bits_mask),
    .io_deq_ready(repeated_repeater_io_deq_ready),
    .io_deq_valid(repeated_repeater_io_deq_valid),
    .io_deq_bits_size(repeated_repeater_io_deq_bits_size),
    .io_deq_bits_source(repeated_repeater_io_deq_bits_source),
    .io_deq_bits_address(repeated_repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeated_repeater_io_deq_bits_mask),
    .io_covSum(repeated_repeater_io_covSum)
  );
  assign auto_in_a_ready = repeated_repeater_io_enq_ready; // @[Nodes.scala 1210:84 Repeater.scala 37:21]
  assign auto_in_d_valid = auto_out_d_valid & last; // @[WidthWidget.scala 71:29]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = {auto_out_d_bits_data,bundleIn_0_d_bits_data_mdata_0}; // @[Cat.scala 31:58]
  assign auto_out_a_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 155:25 156:15]
  assign auto_out_a_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 155:25 156:15]
  assign auto_out_a_bits_source = repeated_repeater_io_deq_bits_source; // @[WidthWidget.scala 155:25 156:15]
  assign auto_out_a_bits_address = repeated_repeater_io_deq_bits_address; // @[WidthWidget.scala 155:25 156:15]
  assign auto_out_a_bits_mask = repeat_sel ? repeat_bundleOut_0_a_bits_mask_mux_1 : repeat_bundleOut_0_a_bits_mask_mux_0
    ; // @[WidthWidget.scala 134:{53,53}]
  assign auto_out_d_ready = auto_in_d_ready | ~last; // @[WidthWidget.scala 70:29]
  assign repeated_repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeated_repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign TLWidthWidget_6_covMap_read_en = 1'h1;
  assign TLWidthWidget_6_covMap_read_addr = TLWidthWidget_6_covState;
  assign TLWidthWidget_6_covMap_read_data = TLWidthWidget_6_covMap[TLWidthWidget_6_covMap_read_addr]; // @[Coverage map for TLWidthWidget_6]
  assign TLWidthWidget_6_covMap_write_data = 1'h1;
  assign TLWidthWidget_6_covMap_write_addr = TLWidthWidget_6_covState;
  assign TLWidthWidget_6_covMap_write_mask = 1'h1;
  assign TLWidthWidget_6_covMap_write_en = ~metaReset;
  assign bundleIn_0_d_bits_data_rdata_written_once_shl = bundleIn_0_d_bits_data_rdata_written_once;
  assign bundleIn_0_d_bits_data_rdata_written_once_pad = {1'h0,bundleIn_0_d_bits_data_rdata_written_once_shl};
  assign count_shl = {count, 1'h0};
  assign count_pad = count_shl;
  assign TLWidthWidget_6_xor0 = bundleIn_0_d_bits_data_rdata_written_once_pad ^ count_pad;
  assign repeated_repeater_sum = TLWidthWidget_6_covSum + repeated_repeater_io_covSum;
  assign io_covSum = repeated_repeater_sum;
  always @(posedge clock) begin
    if (reset) begin // @[WidthWidget.scala 34:27]
      count <= 1'h0; // @[WidthWidget.scala 34:27]
    end else if (_T) begin
      if (last) begin
        count <= 1'h0;
      end else begin
        count <= count + 1'h1;
      end
    end
    if (reset) begin // @[WidthWidget.scala 56:41]
      bundleIn_0_d_bits_data_rdata_written_once <= 1'h0; // @[WidthWidget.scala 56:41]
    end else begin
      bundleIn_0_d_bits_data_rdata_written_once <= _GEN_8;
    end
    if (_T & _bundleOut_0_d_ready_T) begin // @[WidthWidget.scala 63:35]
      if (bundleIn_0_d_bits_data_masked_enable_0) begin
        bundleIn_0_d_bits_data_rdata_0 <= auto_out_d_bits_data;
      end
    end
    TLWidthWidget_6_covState <= TLWidthWidget_6_xor0;
    if (TLWidthWidget_6_covMap_write_en & TLWidthWidget_6_covMap_write_mask) begin
      TLWidthWidget_6_covMap[TLWidthWidget_6_covMap_write_addr] <= TLWidthWidget_6_covMap_write_data; // @[Coverage map for TLWidthWidget_6]
    end
    if (!(TLWidthWidget_6_covMap_read_data | metaReset)) begin
      TLWidthWidget_6_covSum <= TLWidthWidget_6_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    TLWidthWidget_6_covMap[initvar] = 0; //_4[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bundleIn_0_d_bits_data_rdata_written_once = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bundleIn_0_d_bits_data_rdata_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  TLWidthWidget_6_covState = 0; //_3[1:0];
  _RAND_5 = {1{`RANDOM}};
  TLWidthWidget_6_covSum = 0; //_5[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLInterconnectCoupler_11(
  input         clock,
  input         reset,
  input         auto_fragmenter_out_a_ready,
  output        auto_fragmenter_out_a_valid,
  output [1:0]  auto_fragmenter_out_a_bits_size,
  output [11:0] auto_fragmenter_out_a_bits_source,
  output [17:0] auto_fragmenter_out_a_bits_address,
  output        auto_fragmenter_out_d_ready,
  input         auto_fragmenter_out_d_valid,
  input  [1:0]  auto_fragmenter_out_d_bits_size,
  input  [11:0] auto_fragmenter_out_d_bits_source,
  input  [31:0] auto_fragmenter_out_d_bits_data,
  output        auto_tl_in_a_ready,
  input         auto_tl_in_a_valid,
  input  [2:0]  auto_tl_in_a_bits_size,
  input  [6:0]  auto_tl_in_a_bits_source,
  input  [17:0] auto_tl_in_a_bits_address,
  input  [7:0]  auto_tl_in_a_bits_mask,
  input         auto_tl_in_d_ready,
  output        auto_tl_in_d_valid,
  output [2:0]  auto_tl_in_d_bits_size,
  output [6:0]  auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [17:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [3:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [31:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [11:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [17:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [11:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [31:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34]
  wire [29:0] fragmenter_io_covSum; // @[Fragmenter.scala 333:34]
  wire  fragmenter_metaReset; // @[Fragmenter.scala 333:34]
  wire  widget_clock; // @[WidthWidget.scala 219:28]
  wire  widget_reset; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_a_ready; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_a_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_in_a_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_auto_in_a_bits_source; // @[WidthWidget.scala 219:28]
  wire [17:0] widget_auto_in_a_bits_address; // @[WidthWidget.scala 219:28]
  wire [7:0] widget_auto_in_a_bits_mask; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_d_ready; // @[WidthWidget.scala 219:28]
  wire  widget_auto_in_d_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_in_d_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_auto_in_d_bits_source; // @[WidthWidget.scala 219:28]
  wire [63:0] widget_auto_in_d_bits_data; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_a_ready; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_a_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_out_a_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_auto_out_a_bits_source; // @[WidthWidget.scala 219:28]
  wire [17:0] widget_auto_out_a_bits_address; // @[WidthWidget.scala 219:28]
  wire [3:0] widget_auto_out_a_bits_mask; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_d_ready; // @[WidthWidget.scala 219:28]
  wire  widget_auto_out_d_valid; // @[WidthWidget.scala 219:28]
  wire [2:0] widget_auto_out_d_bits_size; // @[WidthWidget.scala 219:28]
  wire [6:0] widget_auto_out_d_bits_source; // @[WidthWidget.scala 219:28]
  wire [31:0] widget_auto_out_d_bits_data; // @[WidthWidget.scala 219:28]
  wire [29:0] widget_io_covSum; // @[WidthWidget.scala 219:28]
  wire  widget_metaReset; // @[WidthWidget.scala 219:28]
  wire [29:0] TLInterconnectCoupler_11_covSum;
  wire [29:0] fragmenter_sum;
  wire [29:0] widget_sum;
  TLFragmenter_4 fragmenter ( // @[Fragmenter.scala 333:34]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .io_covSum(fragmenter_io_covSum),
    .metaReset(fragmenter_metaReset)
  );
  TLWidthWidget_6 widget ( // @[WidthWidget.scala 219:28]
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_size(widget_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_auto_in_d_bits_source),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data),
    .io_covSum(widget_io_covSum),
    .metaReset(widget_metaReset)
  );
  assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_tl_in_a_ready = widget_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_valid = widget_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_size = widget_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_source = widget_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_data = widget_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign fragmenter_clock = clock;
  assign fragmenter_reset = reset;
  assign fragmenter_auto_in_a_valid = widget_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign fragmenter_auto_in_a_bits_size = widget_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fragmenter_auto_in_a_bits_source = widget_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fragmenter_auto_in_a_bits_address = widget_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fragmenter_auto_in_a_bits_mask = widget_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fragmenter_auto_in_d_ready = widget_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign widget_clock = clock;
  assign widget_reset = reset;
  assign widget_auto_in_a_valid = auto_tl_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_size = auto_tl_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_source = auto_tl_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_address = auto_tl_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_mask = auto_tl_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_d_ready = auto_tl_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_ready = fragmenter_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_valid = fragmenter_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_size = fragmenter_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_source = fragmenter_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_data = fragmenter_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign TLInterconnectCoupler_11_covSum = 30'h0;
  assign fragmenter_sum = TLInterconnectCoupler_11_covSum + fragmenter_io_covSum;
  assign widget_sum = fragmenter_sum + widget_io_covSum;
  assign io_covSum = widget_sum;
  assign fragmenter_metaReset = metaReset;
  assign widget_metaReset = metaReset;
endmodule
module Repeater_6(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [6:0]  io_enq_bits_source,
  input  [11:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [6:0]  io_deq_bits_source,
  output [11:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [6:0] saved_source; // @[Repeater.scala 20:18]
  reg [11:0] saved_address; // @[Repeater.scala 20:18]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 19:21 28:{38,45}]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  reg  Repeater_6_covState; // @[Register tracking Repeater_6 state]
  reg  Repeater_6_covMap [0:1]; // @[Coverage map for Repeater_6]
  wire  Repeater_6_covMap_read_en; // @[Coverage map for Repeater_6]
  wire  Repeater_6_covMap_read_addr; // @[Coverage map for Repeater_6]
  wire  Repeater_6_covMap_read_data; // @[Coverage map for Repeater_6]
  wire  Repeater_6_covMap_write_data; // @[Coverage map for Repeater_6]
  wire  Repeater_6_covMap_write_addr; // @[Coverage map for Repeater_6]
  wire  Repeater_6_covMap_write_mask; // @[Coverage map for Repeater_6]
  wire  Repeater_6_covMap_write_en; // @[Coverage map for Repeater_6]
  reg [29:0] Repeater_6_covSum; // @[Sum of coverage map]
  wire  full_shl;
  wire  full_pad;
  assign io_full = full; // @[Repeater.scala 26:11]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21]
  assign Repeater_6_covMap_read_en = 1'h1;
  assign Repeater_6_covMap_read_addr = Repeater_6_covState;
  assign Repeater_6_covMap_read_data = Repeater_6_covMap[Repeater_6_covMap_read_addr]; // @[Coverage map for Repeater_6]
  assign Repeater_6_covMap_write_data = 1'h1;
  assign Repeater_6_covMap_write_addr = Repeater_6_covState;
  assign Repeater_6_covMap_write_mask = 1'h1;
  assign Repeater_6_covMap_write_en = ~metaReset;
  assign full_shl = full;
  assign full_pad = full_shl;
  assign io_covSum = Repeater_6_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin
      full <= 1'h0;
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62]
    end
    Repeater_6_covState <= full_pad;
    if (Repeater_6_covMap_write_en & Repeater_6_covMap_write_mask) begin
      Repeater_6_covMap[Repeater_6_covMap_write_addr] <= Repeater_6_covMap_write_data; // @[Coverage map for Repeater_6]
    end
    if (!(Repeater_6_covMap_read_data | metaReset)) begin
      Repeater_6_covSum <= Repeater_6_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Repeater_6_covMap[initvar] = 0; //_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_source = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  saved_address = _RAND_4[11:0];
  _RAND_5 = {1{`RANDOM}};
  saved_mask = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  Repeater_6_covState = 0; //_6[0:0];
  _RAND_8 = {1{`RANDOM}};
  Repeater_6_covSum = 0; //_8[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_5(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [11:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [1:0]  auto_out_a_bits_size,
  output [10:0] auto_out_a_bits_source,
  output [11:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_size,
  input  [10:0] auto_out_d_bits_source,
  input  [63:0] auto_out_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  repeater_clock; // @[Fragmenter.scala 262:30]
  wire  repeater_reset; // @[Fragmenter.scala 262:30]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_opcode; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30]
  wire [11:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_opcode; // @[Fragmenter.scala 262:30]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30]
  wire [6:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30]
  wire [11:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30]
  wire [7:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30]
  wire [29:0] repeater_io_covSum; // @[Fragmenter.scala 262:30]
  wire  repeater_metaReset; // @[Fragmenter.scala 262:30]
  reg [2:0] acknum; // @[Fragmenter.scala 189:29]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24]
  reg  dToggle; // @[Fragmenter.scala 191:30]
  wire [2:0] dFragnum = auto_out_d_bits_source[2:0]; // @[Fragmenter.scala 192:41]
  wire  dFirst = acknum == 3'h0; // @[Fragmenter.scala 193:29]
  wire  dLast = dFragnum == 3'h0; // @[Fragmenter.scala 194:30]
  wire [3:0] dsizeOH = 4'h1 << auto_out_d_bits_size; // @[OneHot.scala 64:12]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[package.scala 234:46]
  wire  dHasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  _T_5 = ~reset; // @[Fragmenter.scala 202:16]
  wire  ack_decrement = dHasData | dsizeOH[3]; // @[Fragmenter.scala 204:32]
  wire [5:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[Fragmenter.scala 206:47]
  wire [5:0] _GEN_7 = {{3'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69]
  wire [5:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69]
  wire [6:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0}; // @[package.scala 232:35]
  wire [6:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 7'h1; // @[package.scala 232:40]
  wire [6:0] _dFirst_size_T_4 = {1'h0,_dFirst_size_T_1}; // @[Cat.scala 31:58]
  wire [6:0] _dFirst_size_T_5 = ~_dFirst_size_T_4; // @[package.scala 232:53]
  wire [6:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5; // @[package.scala 232:51]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_6[6:4]; // @[OneHot.scala 30:18]
  wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_7 = |dFirst_size_hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28]
  wire [3:0] _dFirst_size_T_8 = _GEN_8 | dFirst_size_lo; // @[OneHot.scala 32:28]
  wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _dFirst_size_T_9 = |dFirst_size_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] dFirst_size = {_dFirst_size_T_7,_dFirst_size_T_9,_dFirst_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  drop = ~dHasData & ~dLast; // @[Fragmenter.scala 222:30]
  wire  bundleOut_0_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35]
  wire  _T_7 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_9 = {{2'd0}, ack_decrement}; // @[Fragmenter.scala 209:55]
  wire [2:0] _acknum_T_1 = acknum - _GEN_9; // @[Fragmenter.scala 209:55]
  wire [2:0] aFrag = repeater_io_deq_bits_size > 3'h3 ? 3'h3 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[package.scala 234:77]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[package.scala 234:46]
  wire  aHasData = ~repeater_io_deq_bits_opcode[2]; // @[Edges.scala 91:28]
  reg [2:0] gennum; // @[Fragmenter.scala 291:29]
  wire  aFirst = gennum == 3'h0; // @[Fragmenter.scala 292:29]
  wire [2:0] _old_gennum1_T_2 = gennum - 3'h1; // @[Fragmenter.scala 293:79]
  wire [2:0] old_gennum1 = aFirst ? aOrigOH1[5:3] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30]
  wire [2:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28]
  wire [2:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26]
  reg  aToggle_r; // @[Reg.scala 16:16]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  aToggle = ~_GEN_5; // @[Fragmenter.scala 297:23]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 50:35]
  wire  _repeater_io_repeat_T = ~aHasData; // @[Fragmenter.scala 302:31]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 3'h0}; // @[Fragmenter.scala 304:65]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88]
  wire [5:0] _GEN_10 = {{3'd0}, aFragOH1}; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10; // @[Fragmenter.scala 304:100]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h7; // @[Fragmenter.scala 304:111]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51]
  wire [11:0] _GEN_11 = {{6'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49]
  wire [7:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,aToggle}; // @[Cat.scala 31:58]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17]
  wire [29:0] TLFragmenter_5_covSum;
  wire [29:0] repeater_sum;
  Repeater_6 repeater ( // @[Fragmenter.scala 262:30]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_opcode(repeater_io_enq_bits_opcode),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_opcode(repeater_io_deq_bits_opcode),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_covSum(repeater_io_covSum),
    .metaReset(repeater_metaReset)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 Fragmenter.scala 263:25]
  assign auto_in_d_valid = auto_out_d_valid & ~drop; // @[Fragmenter.scala 224:36]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32]
  assign auto_in_d_bits_source = auto_out_d_bits_source[10:4]; // @[Fragmenter.scala 226:47]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode; // @[Nodes.scala 1207:84 Fragmenter.scala 303:15]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 Fragmenter.scala 306:25]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 31:58]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11; // @[Fragmenter.scala 304:49]
  assign auto_out_a_bits_mask = repeater_io_full ? 8'hff : auto_in_a_bits_mask; // @[Fragmenter.scala 313:31]
  assign auto_out_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35]
  assign repeater_clock = clock;
  assign repeater_reset = reset;
  assign repeater_io_repeat = ~aHasData & new_gennum != 3'h0; // @[Fragmenter.scala 302:41]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign TLFragmenter_5_covSum = 30'h0;
  assign repeater_sum = TLFragmenter_5_covSum + repeater_io_covSum;
  assign io_covSum = repeater_sum;
  assign repeater_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29]
      acknum <= 3'h0; // @[Fragmenter.scala 189:29]
    end else if (_T_7) begin
      if (dFirst) begin
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29]
      if (dFirst) begin
        dOrig <= dFirst_size;
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30]
    end else if (_T_7) begin
      if (dFirst) begin
        dToggle <= auto_out_d_bits_source[3];
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29]
      gennum <= 3'h0; // @[Fragmenter.scala 291:29]
    end else if (_T_8) begin
      gennum <= new_gennum;
    end
    if (aFirst) begin // @[Reg.scala 17:18]
      aToggle_r <= dToggle; // @[Reg.scala 17:22]
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal; // @[Fragmenter.scala 202:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~repeater_io_full | _repeater_io_repeat_T) & _T_5) begin
          $fatal; // @[Fragmenter.scala 309:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(~repeater_io_full | _repeater_io_repeat_T)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:309 assert (!repeater.io.full || !aHasData)\n"
            ); // @[Fragmenter.scala 309:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_9 | repeater_io_deq_bits_mask == 8'hff) & _T_5) begin
          $fatal; // @[Fragmenter.scala 312:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(_T_9 | repeater_io_deq_bits_mask == 8'hff)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLInterconnectCoupler_12(
  input         clock,
  input         reset,
  input         auto_fragmenter_out_a_ready,
  output        auto_fragmenter_out_a_valid,
  output [2:0]  auto_fragmenter_out_a_bits_opcode,
  output [1:0]  auto_fragmenter_out_a_bits_size,
  output [10:0] auto_fragmenter_out_a_bits_source,
  output [11:0] auto_fragmenter_out_a_bits_address,
  output [7:0]  auto_fragmenter_out_a_bits_mask,
  output        auto_fragmenter_out_d_ready,
  input         auto_fragmenter_out_d_valid,
  input  [2:0]  auto_fragmenter_out_d_bits_opcode,
  input  [1:0]  auto_fragmenter_out_d_bits_size,
  input  [10:0] auto_fragmenter_out_d_bits_source,
  input  [63:0] auto_fragmenter_out_d_bits_data,
  output        auto_tl_in_a_ready,
  input         auto_tl_in_a_valid,
  input  [2:0]  auto_tl_in_a_bits_opcode,
  input  [2:0]  auto_tl_in_a_bits_size,
  input  [6:0]  auto_tl_in_a_bits_source,
  input  [11:0] auto_tl_in_a_bits_address,
  input  [7:0]  auto_tl_in_a_bits_mask,
  input         auto_tl_in_d_ready,
  output        auto_tl_in_d_valid,
  output [2:0]  auto_tl_in_d_bits_opcode,
  output [2:0]  auto_tl_in_d_bits_size,
  output [6:0]  auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [11:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [6:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_out_a_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34]
  wire [11:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34]
  wire [7:0] fragmenter_auto_out_a_bits_mask; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34]
  wire [2:0] fragmenter_auto_out_d_bits_opcode; // @[Fragmenter.scala 333:34]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34]
  wire [10:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34]
  wire [29:0] fragmenter_io_covSum; // @[Fragmenter.scala 333:34]
  wire  fragmenter_metaReset; // @[Fragmenter.scala 333:34]
  wire [29:0] TLInterconnectCoupler_12_covSum;
  wire [29:0] fragmenter_sum;
  TLFragmenter_5 fragmenter ( // @[Fragmenter.scala 333:34]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .io_covSum(fragmenter_io_covSum),
    .metaReset(fragmenter_metaReset)
  );
  assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_opcode = fragmenter_auto_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_a_bits_mask = fragmenter_auto_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_opcode = fragmenter_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign fragmenter_clock = clock;
  assign fragmenter_reset = reset;
  assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_opcode = auto_fragmenter_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign TLInterconnectCoupler_12_covSum = 30'h0;
  assign fragmenter_sum = TLInterconnectCoupler_12_covSum + fragmenter_io_covSum;
  assign io_covSum = fragmenter_sum;
  assign fragmenter_metaReset = metaReset;
endmodule
module PeripheryBus_1(
  input         auto_coupler_to_magic_fragmenter_out_a_ready,
  output        auto_coupler_to_magic_fragmenter_out_a_valid,
  output [2:0]  auto_coupler_to_magic_fragmenter_out_a_bits_opcode,
  output [1:0]  auto_coupler_to_magic_fragmenter_out_a_bits_size,
  output [10:0] auto_coupler_to_magic_fragmenter_out_a_bits_source,
  output [11:0] auto_coupler_to_magic_fragmenter_out_a_bits_address,
  output [7:0]  auto_coupler_to_magic_fragmenter_out_a_bits_mask,
  output        auto_coupler_to_magic_fragmenter_out_d_ready,
  input         auto_coupler_to_magic_fragmenter_out_d_valid,
  input  [2:0]  auto_coupler_to_magic_fragmenter_out_d_bits_opcode,
  input  [1:0]  auto_coupler_to_magic_fragmenter_out_d_bits_size,
  input  [10:0] auto_coupler_to_magic_fragmenter_out_d_bits_source,
  input  [63:0] auto_coupler_to_magic_fragmenter_out_d_bits_data,
  input         auto_coupler_to_MaskROM_fragmenter_out_a_ready,
  output        auto_coupler_to_MaskROM_fragmenter_out_a_valid,
  output [1:0]  auto_coupler_to_MaskROM_fragmenter_out_a_bits_size,
  output [11:0] auto_coupler_to_MaskROM_fragmenter_out_a_bits_source,
  output [17:0] auto_coupler_to_MaskROM_fragmenter_out_a_bits_address,
  output        auto_coupler_to_MaskROM_fragmenter_out_d_ready,
  input         auto_coupler_to_MaskROM_fragmenter_out_d_valid,
  input  [1:0]  auto_coupler_to_MaskROM_fragmenter_out_d_bits_size,
  input  [11:0] auto_coupler_to_MaskROM_fragmenter_out_d_bits_source,
  input  [31:0] auto_coupler_to_MaskROM_fragmenter_out_d_bits_data,
  input         auto_coupler_to_bootrom_fragmenter_out_a_ready,
  output        auto_coupler_to_bootrom_fragmenter_out_a_valid,
  output [1:0]  auto_coupler_to_bootrom_fragmenter_out_a_bits_size,
  output [10:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_source,
  output [16:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_address,
  output        auto_coupler_to_bootrom_fragmenter_out_d_ready,
  input         auto_coupler_to_bootrom_fragmenter_out_d_valid,
  input  [1:0]  auto_coupler_to_bootrom_fragmenter_out_d_bits_size,
  input  [10:0] auto_coupler_to_bootrom_fragmenter_out_d_bits_source,
  input  [63:0] auto_coupler_to_bootrom_fragmenter_out_d_bits_data,
  input         auto_coupler_to_clint_fragmenter_out_a_ready,
  output        auto_coupler_to_clint_fragmenter_out_a_valid,
  output [2:0]  auto_coupler_to_clint_fragmenter_out_a_bits_opcode,
  output [1:0]  auto_coupler_to_clint_fragmenter_out_a_bits_size,
  output [10:0] auto_coupler_to_clint_fragmenter_out_a_bits_source,
  output [25:0] auto_coupler_to_clint_fragmenter_out_a_bits_address,
  output [7:0]  auto_coupler_to_clint_fragmenter_out_a_bits_mask,
  output [63:0] auto_coupler_to_clint_fragmenter_out_a_bits_data,
  output        auto_coupler_to_clint_fragmenter_out_d_ready,
  input         auto_coupler_to_clint_fragmenter_out_d_valid,
  input  [2:0]  auto_coupler_to_clint_fragmenter_out_d_bits_opcode,
  input  [1:0]  auto_coupler_to_clint_fragmenter_out_d_bits_size,
  input  [10:0] auto_coupler_to_clint_fragmenter_out_d_bits_source,
  input  [63:0] auto_coupler_to_clint_fragmenter_out_d_bits_data,
  input         auto_coupler_to_plic_fragmenter_out_a_ready,
  output        auto_coupler_to_plic_fragmenter_out_a_valid,
  output [2:0]  auto_coupler_to_plic_fragmenter_out_a_bits_opcode,
  output [1:0]  auto_coupler_to_plic_fragmenter_out_a_bits_size,
  output [10:0] auto_coupler_to_plic_fragmenter_out_a_bits_source,
  output [27:0] auto_coupler_to_plic_fragmenter_out_a_bits_address,
  output [7:0]  auto_coupler_to_plic_fragmenter_out_a_bits_mask,
  output [63:0] auto_coupler_to_plic_fragmenter_out_a_bits_data,
  output        auto_coupler_to_plic_fragmenter_out_d_ready,
  input         auto_coupler_to_plic_fragmenter_out_d_valid,
  input  [2:0]  auto_coupler_to_plic_fragmenter_out_d_bits_opcode,
  input  [1:0]  auto_coupler_to_plic_fragmenter_out_d_bits_size,
  input  [10:0] auto_coupler_to_plic_fragmenter_out_d_bits_source,
  input  [63:0] auto_coupler_to_plic_fragmenter_out_d_bits_data,
  input         auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready,
  output        auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid,
  output [2:0]  auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode,
  output [2:0]  auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param,
  output [2:0]  auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size,
  output [6:0]  auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source,
  output [30:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address,
  output [7:0]  auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask,
  output [63:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data,
  output        auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready,
  input         auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid,
  input  [2:0]  auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode,
  input  [2:0]  auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size,
  input  [6:0]  auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source,
  input         auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied,
  input  [63:0] auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data,
  input         auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt,
  output        auto_fixedClockNode_out_0_clock,
  output        auto_fixedClockNode_out_0_reset,
  input         auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock,
  input         auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset,
  input         auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock,
  input         auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset,
  output        auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock,
  output        auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset,
  output        auto_bus_xing_in_a_ready,
  input         auto_bus_xing_in_a_valid,
  input  [2:0]  auto_bus_xing_in_a_bits_opcode,
  input  [2:0]  auto_bus_xing_in_a_bits_param,
  input  [3:0]  auto_bus_xing_in_a_bits_size,
  input  [6:0]  auto_bus_xing_in_a_bits_source,
  input  [30:0] auto_bus_xing_in_a_bits_address,
  input  [7:0]  auto_bus_xing_in_a_bits_mask,
  input  [63:0] auto_bus_xing_in_a_bits_data,
  input         auto_bus_xing_in_d_ready,
  output        auto_bus_xing_in_d_valid,
  output [2:0]  auto_bus_xing_in_d_bits_opcode,
  output [3:0]  auto_bus_xing_in_d_bits_size,
  output [6:0]  auto_bus_xing_in_d_bits_source,
  output        auto_bus_xing_in_d_bits_denied,
  output [63:0] auto_bus_xing_in_d_bits_data,
  output        auto_bus_xing_in_d_bits_corrupt,
  output        clock,
  output        reset,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_clock;
  wire  subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_reset;
  wire  subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_clock;
  wire  subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_reset;
  wire  subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_clock;
  wire  subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_reset;
  wire  subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_clock;
  wire  subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_reset;
  wire  clockGroup_auto_in_member_subsystem_cbus_0_clock;
  wire  clockGroup_auto_in_member_subsystem_cbus_0_reset;
  wire  clockGroup_auto_out_clock;
  wire  clockGroup_auto_out_reset;
  wire  fixedClockNode_auto_in_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_in_reset; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_2_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_2_reset; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_1_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_1_reset; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_0_clock; // @[ClockGroup.scala 106:107]
  wire  fixedClockNode_auto_out_0_reset; // @[ClockGroup.scala 106:107]
  wire [29:0] fixedClockNode_io_covSum; // @[ClockGroup.scala 106:107]
  wire  fixer_clock; // @[PeripheryBus.scala 47:33]
  wire  fixer_reset; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_in_a_ready; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_in_a_valid; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_in_a_bits_opcode; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_in_a_bits_param; // @[PeripheryBus.scala 47:33]
  wire [3:0] fixer_auto_in_a_bits_size; // @[PeripheryBus.scala 47:33]
  wire [6:0] fixer_auto_in_a_bits_source; // @[PeripheryBus.scala 47:33]
  wire [30:0] fixer_auto_in_a_bits_address; // @[PeripheryBus.scala 47:33]
  wire [7:0] fixer_auto_in_a_bits_mask; // @[PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_in_a_bits_data; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_in_d_ready; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_in_d_valid; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_in_d_bits_opcode; // @[PeripheryBus.scala 47:33]
  wire [3:0] fixer_auto_in_d_bits_size; // @[PeripheryBus.scala 47:33]
  wire [6:0] fixer_auto_in_d_bits_source; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_in_d_bits_denied; // @[PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_in_d_bits_data; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_in_d_bits_corrupt; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_a_ready; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_a_valid; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_out_a_bits_opcode; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_out_a_bits_param; // @[PeripheryBus.scala 47:33]
  wire [3:0] fixer_auto_out_a_bits_size; // @[PeripheryBus.scala 47:33]
  wire [6:0] fixer_auto_out_a_bits_source; // @[PeripheryBus.scala 47:33]
  wire [30:0] fixer_auto_out_a_bits_address; // @[PeripheryBus.scala 47:33]
  wire [7:0] fixer_auto_out_a_bits_mask; // @[PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_out_a_bits_data; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_d_ready; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_d_valid; // @[PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_out_d_bits_opcode; // @[PeripheryBus.scala 47:33]
  wire [3:0] fixer_auto_out_d_bits_size; // @[PeripheryBus.scala 47:33]
  wire [6:0] fixer_auto_out_d_bits_source; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_d_bits_denied; // @[PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_out_d_bits_data; // @[PeripheryBus.scala 47:33]
  wire  fixer_auto_out_d_bits_corrupt; // @[PeripheryBus.scala 47:33]
  wire [29:0] fixer_io_covSum; // @[PeripheryBus.scala 47:33]
  wire  fixer_metaReset; // @[PeripheryBus.scala 47:33]
  wire  in_xbar_auto_in_a_ready;
  wire  in_xbar_auto_in_a_valid;
  wire [2:0] in_xbar_auto_in_a_bits_opcode;
  wire [2:0] in_xbar_auto_in_a_bits_param;
  wire [3:0] in_xbar_auto_in_a_bits_size;
  wire [6:0] in_xbar_auto_in_a_bits_source;
  wire [30:0] in_xbar_auto_in_a_bits_address;
  wire [7:0] in_xbar_auto_in_a_bits_mask;
  wire [63:0] in_xbar_auto_in_a_bits_data;
  wire  in_xbar_auto_in_d_ready;
  wire  in_xbar_auto_in_d_valid;
  wire [2:0] in_xbar_auto_in_d_bits_opcode;
  wire [3:0] in_xbar_auto_in_d_bits_size;
  wire [6:0] in_xbar_auto_in_d_bits_source;
  wire  in_xbar_auto_in_d_bits_denied;
  wire [63:0] in_xbar_auto_in_d_bits_data;
  wire  in_xbar_auto_in_d_bits_corrupt;
  wire  in_xbar_auto_out_a_ready;
  wire  in_xbar_auto_out_a_valid;
  wire [2:0] in_xbar_auto_out_a_bits_opcode;
  wire [2:0] in_xbar_auto_out_a_bits_param;
  wire [3:0] in_xbar_auto_out_a_bits_size;
  wire [6:0] in_xbar_auto_out_a_bits_source;
  wire [30:0] in_xbar_auto_out_a_bits_address;
  wire [7:0] in_xbar_auto_out_a_bits_mask;
  wire [63:0] in_xbar_auto_out_a_bits_data;
  wire  in_xbar_auto_out_d_ready;
  wire  in_xbar_auto_out_d_valid;
  wire [2:0] in_xbar_auto_out_d_bits_opcode;
  wire [3:0] in_xbar_auto_out_d_bits_size;
  wire [6:0] in_xbar_auto_out_d_bits_source;
  wire  in_xbar_auto_out_d_bits_denied;
  wire [63:0] in_xbar_auto_out_d_bits_data;
  wire  in_xbar_auto_out_d_bits_corrupt;
  wire  out_xbar_clock; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_reset; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_a_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_a_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_in_a_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_in_a_bits_param; // @[PeripheryBus.scala 50:30]
  wire [3:0] out_xbar_auto_in_a_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_in_a_bits_source; // @[PeripheryBus.scala 50:30]
  wire [30:0] out_xbar_auto_in_a_bits_address; // @[PeripheryBus.scala 50:30]
  wire [7:0] out_xbar_auto_in_a_bits_mask; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_in_a_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_d_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_d_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_in_d_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [3:0] out_xbar_auto_in_d_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_in_d_bits_source; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_d_bits_denied; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_in_d_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_d_bits_corrupt; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_6_a_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_6_a_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_6_a_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_6_a_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_6_a_bits_source; // @[PeripheryBus.scala 50:30]
  wire [11:0] out_xbar_auto_out_6_a_bits_address; // @[PeripheryBus.scala 50:30]
  wire [7:0] out_xbar_auto_out_6_a_bits_mask; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_6_d_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_6_d_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_6_d_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_6_d_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_6_d_bits_source; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_6_d_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_5_a_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_5_a_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_5_a_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_5_a_bits_source; // @[PeripheryBus.scala 50:30]
  wire [17:0] out_xbar_auto_out_5_a_bits_address; // @[PeripheryBus.scala 50:30]
  wire [7:0] out_xbar_auto_out_5_a_bits_mask; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_5_d_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_5_d_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_5_d_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_5_d_bits_source; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_5_d_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_4_a_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_4_a_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_4_a_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_4_a_bits_source; // @[PeripheryBus.scala 50:30]
  wire [16:0] out_xbar_auto_out_4_a_bits_address; // @[PeripheryBus.scala 50:30]
  wire [7:0] out_xbar_auto_out_4_a_bits_mask; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_4_d_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_4_d_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_4_d_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_4_d_bits_source; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_4_d_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_3_a_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_3_a_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_3_a_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_3_a_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_3_a_bits_source; // @[PeripheryBus.scala 50:30]
  wire [25:0] out_xbar_auto_out_3_a_bits_address; // @[PeripheryBus.scala 50:30]
  wire [7:0] out_xbar_auto_out_3_a_bits_mask; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_3_a_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_3_d_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_3_d_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_3_d_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_3_d_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_3_d_bits_source; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_3_d_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_2_a_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_2_a_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_2_a_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_2_a_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_2_a_bits_source; // @[PeripheryBus.scala 50:30]
  wire [27:0] out_xbar_auto_out_2_a_bits_address; // @[PeripheryBus.scala 50:30]
  wire [7:0] out_xbar_auto_out_2_a_bits_mask; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_2_a_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_2_d_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_2_d_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_2_d_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_2_d_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_2_d_bits_source; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_2_d_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_1_a_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_1_a_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_1_a_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_1_a_bits_param; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_1_a_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_1_a_bits_source; // @[PeripheryBus.scala 50:30]
  wire [30:0] out_xbar_auto_out_1_a_bits_address; // @[PeripheryBus.scala 50:30]
  wire [7:0] out_xbar_auto_out_1_a_bits_mask; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_1_a_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_1_d_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_1_d_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_1_d_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_1_d_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_1_d_bits_source; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_1_d_bits_denied; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_1_d_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_1_d_bits_corrupt; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_0_a_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_0_a_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_0_a_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [3:0] out_xbar_auto_out_0_a_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_0_a_bits_source; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_0_d_ready; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_0_d_valid; // @[PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_0_d_bits_opcode; // @[PeripheryBus.scala 50:30]
  wire [3:0] out_xbar_auto_out_0_d_bits_size; // @[PeripheryBus.scala 50:30]
  wire [6:0] out_xbar_auto_out_0_d_bits_source; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_0_d_bits_denied; // @[PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_0_d_bits_data; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_0_d_bits_corrupt; // @[PeripheryBus.scala 50:30]
  wire [29:0] out_xbar_io_covSum; // @[PeripheryBus.scala 50:30]
  wire  out_xbar_metaReset; // @[PeripheryBus.scala 50:30]
  wire  buffer_clock; // @[Buffer.scala 68:28]
  wire  buffer_reset; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28]
  wire [30:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28]
  wire [30:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28]
  wire [6:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire [29:0] buffer_io_covSum; // @[Buffer.scala 68:28]
  wire  atomics_clock; // @[AtomicAutomata.scala 283:29]
  wire  atomics_reset; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_a_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_a_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_a_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_a_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [3:0] atomics_auto_in_a_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_in_a_bits_source; // @[AtomicAutomata.scala 283:29]
  wire [30:0] atomics_auto_in_a_bits_address; // @[AtomicAutomata.scala 283:29]
  wire [7:0] atomics_auto_in_a_bits_mask; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_in_a_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_in_d_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [3:0] atomics_auto_in_d_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_in_d_bits_source; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_bits_denied; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_in_d_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_in_d_bits_corrupt; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_a_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_a_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_a_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_a_bits_param; // @[AtomicAutomata.scala 283:29]
  wire [3:0] atomics_auto_out_a_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_out_a_bits_source; // @[AtomicAutomata.scala 283:29]
  wire [30:0] atomics_auto_out_a_bits_address; // @[AtomicAutomata.scala 283:29]
  wire [7:0] atomics_auto_out_a_bits_mask; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_out_a_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_ready; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_valid; // @[AtomicAutomata.scala 283:29]
  wire [2:0] atomics_auto_out_d_bits_opcode; // @[AtomicAutomata.scala 283:29]
  wire [3:0] atomics_auto_out_d_bits_size; // @[AtomicAutomata.scala 283:29]
  wire [6:0] atomics_auto_out_d_bits_source; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_bits_denied; // @[AtomicAutomata.scala 283:29]
  wire [63:0] atomics_auto_out_d_bits_data; // @[AtomicAutomata.scala 283:29]
  wire  atomics_auto_out_d_bits_corrupt; // @[AtomicAutomata.scala 283:29]
  wire [29:0] atomics_io_covSum; // @[AtomicAutomata.scala 283:29]
  wire  atomics_metaReset; // @[AtomicAutomata.scala 283:29]
  wire  wrapped_error_device_clock; // @[LazyModule.scala 432:27]
  wire  wrapped_error_device_reset; // @[LazyModule.scala 432:27]
  wire  wrapped_error_device_auto_buffer_in_a_ready; // @[LazyModule.scala 432:27]
  wire  wrapped_error_device_auto_buffer_in_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] wrapped_error_device_auto_buffer_in_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [3:0] wrapped_error_device_auto_buffer_in_a_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] wrapped_error_device_auto_buffer_in_a_bits_source; // @[LazyModule.scala 432:27]
  wire  wrapped_error_device_auto_buffer_in_d_ready; // @[LazyModule.scala 432:27]
  wire  wrapped_error_device_auto_buffer_in_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] wrapped_error_device_auto_buffer_in_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [3:0] wrapped_error_device_auto_buffer_in_d_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] wrapped_error_device_auto_buffer_in_d_bits_source; // @[LazyModule.scala 432:27]
  wire  wrapped_error_device_auto_buffer_in_d_bits_denied; // @[LazyModule.scala 432:27]
  wire [63:0] wrapped_error_device_auto_buffer_in_d_bits_data; // @[LazyModule.scala 432:27]
  wire  wrapped_error_device_auto_buffer_in_d_bits_corrupt; // @[LazyModule.scala 432:27]
  wire [29:0] wrapped_error_device_io_covSum; // @[LazyModule.scala 432:27]
  wire  buffer_1_auto_in_a_ready;
  wire  buffer_1_auto_in_a_valid;
  wire [2:0] buffer_1_auto_in_a_bits_opcode;
  wire [2:0] buffer_1_auto_in_a_bits_param;
  wire [3:0] buffer_1_auto_in_a_bits_size;
  wire [6:0] buffer_1_auto_in_a_bits_source;
  wire [30:0] buffer_1_auto_in_a_bits_address;
  wire [7:0] buffer_1_auto_in_a_bits_mask;
  wire [63:0] buffer_1_auto_in_a_bits_data;
  wire  buffer_1_auto_in_d_ready;
  wire  buffer_1_auto_in_d_valid;
  wire [2:0] buffer_1_auto_in_d_bits_opcode;
  wire [3:0] buffer_1_auto_in_d_bits_size;
  wire [6:0] buffer_1_auto_in_d_bits_source;
  wire  buffer_1_auto_in_d_bits_denied;
  wire [63:0] buffer_1_auto_in_d_bits_data;
  wire  buffer_1_auto_in_d_bits_corrupt;
  wire  buffer_1_auto_out_a_ready;
  wire  buffer_1_auto_out_a_valid;
  wire [2:0] buffer_1_auto_out_a_bits_opcode;
  wire [2:0] buffer_1_auto_out_a_bits_param;
  wire [3:0] buffer_1_auto_out_a_bits_size;
  wire [6:0] buffer_1_auto_out_a_bits_source;
  wire [30:0] buffer_1_auto_out_a_bits_address;
  wire [7:0] buffer_1_auto_out_a_bits_mask;
  wire [63:0] buffer_1_auto_out_a_bits_data;
  wire  buffer_1_auto_out_d_ready;
  wire  buffer_1_auto_out_d_valid;
  wire [2:0] buffer_1_auto_out_d_bits_opcode;
  wire [3:0] buffer_1_auto_out_d_bits_size;
  wire [6:0] buffer_1_auto_out_d_bits_source;
  wire  buffer_1_auto_out_d_bits_denied;
  wire [63:0] buffer_1_auto_out_d_bits_data;
  wire  buffer_1_auto_out_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_ready;
  wire  coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_param;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_source;
  wire [30:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_address;
  wire [7:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_data;
  wire  coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_ready;
  wire  coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_source;
  wire  coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_data;
  wire  coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_ready;
  wire  coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_param;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_source;
  wire [30:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_address;
  wire [7:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_data;
  wire  coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_ready;
  wire  coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_source;
  wire  coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_data;
  wire  coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_ready;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_param;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_source;
  wire [30:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_address;
  wire [7:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_data;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_ready;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_source;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_data;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_ready;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_param;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_source;
  wire [30:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_address;
  wire [7:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_data;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_ready;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_size;
  wire [6:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_source;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_data;
  wire  coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_corrupt;
  wire  coupler_to_plic_clock; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_reset; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_auto_fragmenter_out_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_auto_fragmenter_out_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_plic_auto_fragmenter_out_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_plic_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_plic_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 432:27]
  wire [27:0] coupler_to_plic_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_plic_auto_fragmenter_out_a_bits_mask; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_plic_auto_fragmenter_out_a_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_auto_fragmenter_out_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_auto_fragmenter_out_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_plic_auto_fragmenter_out_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_plic_auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_plic_auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_plic_auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_auto_tl_in_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_auto_tl_in_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_plic_auto_tl_in_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_plic_auto_tl_in_a_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_plic_auto_tl_in_a_bits_source; // @[LazyModule.scala 432:27]
  wire [27:0] coupler_to_plic_auto_tl_in_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_plic_auto_tl_in_a_bits_mask; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_plic_auto_tl_in_a_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_auto_tl_in_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_auto_tl_in_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_plic_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_plic_auto_tl_in_d_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_plic_auto_tl_in_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_plic_auto_tl_in_d_bits_data; // @[LazyModule.scala 432:27]
  wire [29:0] coupler_to_plic_io_covSum; // @[LazyModule.scala 432:27]
  wire  coupler_to_plic_metaReset; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_clock; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_reset; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_auto_fragmenter_out_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_auto_fragmenter_out_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_clint_auto_fragmenter_out_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_clint_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_clint_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 432:27]
  wire [25:0] coupler_to_clint_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_clint_auto_fragmenter_out_a_bits_mask; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_clint_auto_fragmenter_out_a_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_auto_fragmenter_out_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_auto_fragmenter_out_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_clint_auto_fragmenter_out_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_clint_auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_clint_auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_clint_auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_auto_tl_in_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_auto_tl_in_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_clint_auto_tl_in_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_clint_auto_tl_in_a_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_clint_auto_tl_in_a_bits_source; // @[LazyModule.scala 432:27]
  wire [25:0] coupler_to_clint_auto_tl_in_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_clint_auto_tl_in_a_bits_mask; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_clint_auto_tl_in_a_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_auto_tl_in_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_auto_tl_in_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_clint_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_clint_auto_tl_in_d_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_clint_auto_tl_in_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_clint_auto_tl_in_d_bits_data; // @[LazyModule.scala 432:27]
  wire [29:0] coupler_to_clint_io_covSum; // @[LazyModule.scala 432:27]
  wire  coupler_to_clint_metaReset; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_clock; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_reset; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_auto_fragmenter_out_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_auto_fragmenter_out_a_valid; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 432:27]
  wire [16:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_auto_fragmenter_out_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_auto_fragmenter_out_d_valid; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_bootrom_auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_bootrom_auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_bootrom_auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_auto_tl_in_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_auto_tl_in_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_bootrom_auto_tl_in_a_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_bootrom_auto_tl_in_a_bits_source; // @[LazyModule.scala 432:27]
  wire [16:0] coupler_to_bootrom_auto_tl_in_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_bootrom_auto_tl_in_a_bits_mask; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_auto_tl_in_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_auto_tl_in_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_bootrom_auto_tl_in_d_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_bootrom_auto_tl_in_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_bootrom_auto_tl_in_d_bits_data; // @[LazyModule.scala 432:27]
  wire [29:0] coupler_to_bootrom_io_covSum; // @[LazyModule.scala 432:27]
  wire  coupler_to_bootrom_metaReset; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_clock; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_reset; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_auto_fragmenter_out_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_auto_fragmenter_out_a_valid; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_MaskROM_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 432:27]
  wire [11:0] coupler_to_MaskROM_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 432:27]
  wire [17:0] coupler_to_MaskROM_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_auto_fragmenter_out_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_auto_fragmenter_out_d_valid; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_MaskROM_auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 432:27]
  wire [11:0] coupler_to_MaskROM_auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 432:27]
  wire [31:0] coupler_to_MaskROM_auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_auto_tl_in_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_auto_tl_in_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_MaskROM_auto_tl_in_a_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_MaskROM_auto_tl_in_a_bits_source; // @[LazyModule.scala 432:27]
  wire [17:0] coupler_to_MaskROM_auto_tl_in_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_MaskROM_auto_tl_in_a_bits_mask; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_auto_tl_in_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_auto_tl_in_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_MaskROM_auto_tl_in_d_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_MaskROM_auto_tl_in_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_MaskROM_auto_tl_in_d_bits_data; // @[LazyModule.scala 432:27]
  wire [29:0] coupler_to_MaskROM_io_covSum; // @[LazyModule.scala 432:27]
  wire  coupler_to_MaskROM_metaReset; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_clock; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_reset; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_auto_fragmenter_out_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_auto_fragmenter_out_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_magic_auto_fragmenter_out_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_magic_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_magic_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 432:27]
  wire [11:0] coupler_to_magic_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_magic_auto_fragmenter_out_a_bits_mask; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_auto_fragmenter_out_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_auto_fragmenter_out_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_magic_auto_fragmenter_out_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_magic_auto_fragmenter_out_d_bits_size; // @[LazyModule.scala 432:27]
  wire [10:0] coupler_to_magic_auto_fragmenter_out_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_magic_auto_fragmenter_out_d_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_auto_tl_in_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_auto_tl_in_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_magic_auto_tl_in_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_magic_auto_tl_in_a_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_magic_auto_tl_in_a_bits_source; // @[LazyModule.scala 432:27]
  wire [11:0] coupler_to_magic_auto_tl_in_a_bits_address; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_magic_auto_tl_in_a_bits_mask; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_auto_tl_in_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_auto_tl_in_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_magic_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_magic_auto_tl_in_d_bits_size; // @[LazyModule.scala 432:27]
  wire [6:0] coupler_to_magic_auto_tl_in_d_bits_source; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_magic_auto_tl_in_d_bits_data; // @[LazyModule.scala 432:27]
  wire [29:0] coupler_to_magic_io_covSum; // @[LazyModule.scala 432:27]
  wire  coupler_to_magic_metaReset; // @[LazyModule.scala 432:27]
  wire [29:0] PeripheryBus_1_covSum;
  wire [29:0] atomics_sum;
  wire [29:0] coupler_to_clint_sum;
  wire [29:0] wrapped_error_device_sum;
  wire [29:0] fixedClockNode_sum;
  wire [29:0] fixer_sum;
  wire [29:0] coupler_to_bootrom_sum;
  wire [29:0] out_xbar_sum;
  wire [29:0] coupler_to_magic_sum;
  wire [29:0] coupler_to_plic_sum;
  wire [29:0] coupler_to_MaskROM_sum;
  wire [29:0] buffer_sum;
  FixedClockBroadcast fixedClockNode ( // @[ClockGroup.scala 106:107]
    .auto_in_clock(fixedClockNode_auto_in_clock),
    .auto_in_reset(fixedClockNode_auto_in_reset),
    .auto_out_2_clock(fixedClockNode_auto_out_2_clock),
    .auto_out_2_reset(fixedClockNode_auto_out_2_reset),
    .auto_out_1_clock(fixedClockNode_auto_out_1_clock),
    .auto_out_1_reset(fixedClockNode_auto_out_1_reset),
    .auto_out_0_clock(fixedClockNode_auto_out_0_clock),
    .auto_out_0_reset(fixedClockNode_auto_out_0_reset),
    .io_covSum(fixedClockNode_io_covSum)
  );
  TLFIFOFixer_3 fixer ( // @[PeripheryBus.scala 47:33]
    .clock(fixer_clock),
    .reset(fixer_reset),
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fixer_auto_in_a_bits_param),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_auto_in_a_bits_data),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fixer_auto_out_a_bits_param),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_auto_out_a_bits_data),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt),
    .io_covSum(fixer_io_covSum),
    .metaReset(fixer_metaReset)
  );
  TLXbar_5 out_xbar ( // @[PeripheryBus.scala 50:30]
    .clock(out_xbar_clock),
    .reset(out_xbar_reset),
    .auto_in_a_ready(out_xbar_auto_in_a_ready),
    .auto_in_a_valid(out_xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(out_xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(out_xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(out_xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(out_xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(out_xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(out_xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(out_xbar_auto_in_a_bits_data),
    .auto_in_d_ready(out_xbar_auto_in_d_ready),
    .auto_in_d_valid(out_xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(out_xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(out_xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(out_xbar_auto_in_d_bits_source),
    .auto_in_d_bits_denied(out_xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(out_xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(out_xbar_auto_in_d_bits_corrupt),
    .auto_out_6_a_ready(out_xbar_auto_out_6_a_ready),
    .auto_out_6_a_valid(out_xbar_auto_out_6_a_valid),
    .auto_out_6_a_bits_opcode(out_xbar_auto_out_6_a_bits_opcode),
    .auto_out_6_a_bits_size(out_xbar_auto_out_6_a_bits_size),
    .auto_out_6_a_bits_source(out_xbar_auto_out_6_a_bits_source),
    .auto_out_6_a_bits_address(out_xbar_auto_out_6_a_bits_address),
    .auto_out_6_a_bits_mask(out_xbar_auto_out_6_a_bits_mask),
    .auto_out_6_d_ready(out_xbar_auto_out_6_d_ready),
    .auto_out_6_d_valid(out_xbar_auto_out_6_d_valid),
    .auto_out_6_d_bits_opcode(out_xbar_auto_out_6_d_bits_opcode),
    .auto_out_6_d_bits_size(out_xbar_auto_out_6_d_bits_size),
    .auto_out_6_d_bits_source(out_xbar_auto_out_6_d_bits_source),
    .auto_out_6_d_bits_data(out_xbar_auto_out_6_d_bits_data),
    .auto_out_5_a_ready(out_xbar_auto_out_5_a_ready),
    .auto_out_5_a_valid(out_xbar_auto_out_5_a_valid),
    .auto_out_5_a_bits_size(out_xbar_auto_out_5_a_bits_size),
    .auto_out_5_a_bits_source(out_xbar_auto_out_5_a_bits_source),
    .auto_out_5_a_bits_address(out_xbar_auto_out_5_a_bits_address),
    .auto_out_5_a_bits_mask(out_xbar_auto_out_5_a_bits_mask),
    .auto_out_5_d_ready(out_xbar_auto_out_5_d_ready),
    .auto_out_5_d_valid(out_xbar_auto_out_5_d_valid),
    .auto_out_5_d_bits_size(out_xbar_auto_out_5_d_bits_size),
    .auto_out_5_d_bits_source(out_xbar_auto_out_5_d_bits_source),
    .auto_out_5_d_bits_data(out_xbar_auto_out_5_d_bits_data),
    .auto_out_4_a_ready(out_xbar_auto_out_4_a_ready),
    .auto_out_4_a_valid(out_xbar_auto_out_4_a_valid),
    .auto_out_4_a_bits_size(out_xbar_auto_out_4_a_bits_size),
    .auto_out_4_a_bits_source(out_xbar_auto_out_4_a_bits_source),
    .auto_out_4_a_bits_address(out_xbar_auto_out_4_a_bits_address),
    .auto_out_4_a_bits_mask(out_xbar_auto_out_4_a_bits_mask),
    .auto_out_4_d_ready(out_xbar_auto_out_4_d_ready),
    .auto_out_4_d_valid(out_xbar_auto_out_4_d_valid),
    .auto_out_4_d_bits_size(out_xbar_auto_out_4_d_bits_size),
    .auto_out_4_d_bits_source(out_xbar_auto_out_4_d_bits_source),
    .auto_out_4_d_bits_data(out_xbar_auto_out_4_d_bits_data),
    .auto_out_3_a_ready(out_xbar_auto_out_3_a_ready),
    .auto_out_3_a_valid(out_xbar_auto_out_3_a_valid),
    .auto_out_3_a_bits_opcode(out_xbar_auto_out_3_a_bits_opcode),
    .auto_out_3_a_bits_size(out_xbar_auto_out_3_a_bits_size),
    .auto_out_3_a_bits_source(out_xbar_auto_out_3_a_bits_source),
    .auto_out_3_a_bits_address(out_xbar_auto_out_3_a_bits_address),
    .auto_out_3_a_bits_mask(out_xbar_auto_out_3_a_bits_mask),
    .auto_out_3_a_bits_data(out_xbar_auto_out_3_a_bits_data),
    .auto_out_3_d_ready(out_xbar_auto_out_3_d_ready),
    .auto_out_3_d_valid(out_xbar_auto_out_3_d_valid),
    .auto_out_3_d_bits_opcode(out_xbar_auto_out_3_d_bits_opcode),
    .auto_out_3_d_bits_size(out_xbar_auto_out_3_d_bits_size),
    .auto_out_3_d_bits_source(out_xbar_auto_out_3_d_bits_source),
    .auto_out_3_d_bits_data(out_xbar_auto_out_3_d_bits_data),
    .auto_out_2_a_ready(out_xbar_auto_out_2_a_ready),
    .auto_out_2_a_valid(out_xbar_auto_out_2_a_valid),
    .auto_out_2_a_bits_opcode(out_xbar_auto_out_2_a_bits_opcode),
    .auto_out_2_a_bits_size(out_xbar_auto_out_2_a_bits_size),
    .auto_out_2_a_bits_source(out_xbar_auto_out_2_a_bits_source),
    .auto_out_2_a_bits_address(out_xbar_auto_out_2_a_bits_address),
    .auto_out_2_a_bits_mask(out_xbar_auto_out_2_a_bits_mask),
    .auto_out_2_a_bits_data(out_xbar_auto_out_2_a_bits_data),
    .auto_out_2_d_ready(out_xbar_auto_out_2_d_ready),
    .auto_out_2_d_valid(out_xbar_auto_out_2_d_valid),
    .auto_out_2_d_bits_opcode(out_xbar_auto_out_2_d_bits_opcode),
    .auto_out_2_d_bits_size(out_xbar_auto_out_2_d_bits_size),
    .auto_out_2_d_bits_source(out_xbar_auto_out_2_d_bits_source),
    .auto_out_2_d_bits_data(out_xbar_auto_out_2_d_bits_data),
    .auto_out_1_a_ready(out_xbar_auto_out_1_a_ready),
    .auto_out_1_a_valid(out_xbar_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(out_xbar_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_param(out_xbar_auto_out_1_a_bits_param),
    .auto_out_1_a_bits_size(out_xbar_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(out_xbar_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(out_xbar_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_mask(out_xbar_auto_out_1_a_bits_mask),
    .auto_out_1_a_bits_data(out_xbar_auto_out_1_a_bits_data),
    .auto_out_1_d_ready(out_xbar_auto_out_1_d_ready),
    .auto_out_1_d_valid(out_xbar_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(out_xbar_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_size(out_xbar_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(out_xbar_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_denied(out_xbar_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_data(out_xbar_auto_out_1_d_bits_data),
    .auto_out_1_d_bits_corrupt(out_xbar_auto_out_1_d_bits_corrupt),
    .auto_out_0_a_ready(out_xbar_auto_out_0_a_ready),
    .auto_out_0_a_valid(out_xbar_auto_out_0_a_valid),
    .auto_out_0_a_bits_opcode(out_xbar_auto_out_0_a_bits_opcode),
    .auto_out_0_a_bits_size(out_xbar_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(out_xbar_auto_out_0_a_bits_source),
    .auto_out_0_d_ready(out_xbar_auto_out_0_d_ready),
    .auto_out_0_d_valid(out_xbar_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(out_xbar_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_size(out_xbar_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(out_xbar_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_denied(out_xbar_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_data(out_xbar_auto_out_0_d_bits_data),
    .auto_out_0_d_bits_corrupt(out_xbar_auto_out_0_d_bits_corrupt),
    .io_covSum(out_xbar_io_covSum),
    .metaReset(out_xbar_metaReset)
  );
  TLBuffer_4 buffer ( // @[Buffer.scala 68:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt),
    .io_covSum(buffer_io_covSum)
  );
  TLAtomicAutomata_1 atomics ( // @[AtomicAutomata.scala 283:29]
    .clock(atomics_clock),
    .reset(atomics_reset),
    .auto_in_a_ready(atomics_auto_in_a_ready),
    .auto_in_a_valid(atomics_auto_in_a_valid),
    .auto_in_a_bits_opcode(atomics_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(atomics_auto_in_a_bits_param),
    .auto_in_a_bits_size(atomics_auto_in_a_bits_size),
    .auto_in_a_bits_source(atomics_auto_in_a_bits_source),
    .auto_in_a_bits_address(atomics_auto_in_a_bits_address),
    .auto_in_a_bits_mask(atomics_auto_in_a_bits_mask),
    .auto_in_a_bits_data(atomics_auto_in_a_bits_data),
    .auto_in_d_ready(atomics_auto_in_d_ready),
    .auto_in_d_valid(atomics_auto_in_d_valid),
    .auto_in_d_bits_opcode(atomics_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(atomics_auto_in_d_bits_size),
    .auto_in_d_bits_source(atomics_auto_in_d_bits_source),
    .auto_in_d_bits_denied(atomics_auto_in_d_bits_denied),
    .auto_in_d_bits_data(atomics_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(atomics_auto_in_d_bits_corrupt),
    .auto_out_a_ready(atomics_auto_out_a_ready),
    .auto_out_a_valid(atomics_auto_out_a_valid),
    .auto_out_a_bits_opcode(atomics_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(atomics_auto_out_a_bits_param),
    .auto_out_a_bits_size(atomics_auto_out_a_bits_size),
    .auto_out_a_bits_source(atomics_auto_out_a_bits_source),
    .auto_out_a_bits_address(atomics_auto_out_a_bits_address),
    .auto_out_a_bits_mask(atomics_auto_out_a_bits_mask),
    .auto_out_a_bits_data(atomics_auto_out_a_bits_data),
    .auto_out_d_ready(atomics_auto_out_d_ready),
    .auto_out_d_valid(atomics_auto_out_d_valid),
    .auto_out_d_bits_opcode(atomics_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(atomics_auto_out_d_bits_size),
    .auto_out_d_bits_source(atomics_auto_out_d_bits_source),
    .auto_out_d_bits_denied(atomics_auto_out_d_bits_denied),
    .auto_out_d_bits_data(atomics_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(atomics_auto_out_d_bits_corrupt),
    .io_covSum(atomics_io_covSum),
    .metaReset(atomics_metaReset)
  );
  ErrorDeviceWrapper wrapped_error_device ( // @[LazyModule.scala 432:27]
    .clock(wrapped_error_device_clock),
    .reset(wrapped_error_device_reset),
    .auto_buffer_in_a_ready(wrapped_error_device_auto_buffer_in_a_ready),
    .auto_buffer_in_a_valid(wrapped_error_device_auto_buffer_in_a_valid),
    .auto_buffer_in_a_bits_opcode(wrapped_error_device_auto_buffer_in_a_bits_opcode),
    .auto_buffer_in_a_bits_size(wrapped_error_device_auto_buffer_in_a_bits_size),
    .auto_buffer_in_a_bits_source(wrapped_error_device_auto_buffer_in_a_bits_source),
    .auto_buffer_in_d_ready(wrapped_error_device_auto_buffer_in_d_ready),
    .auto_buffer_in_d_valid(wrapped_error_device_auto_buffer_in_d_valid),
    .auto_buffer_in_d_bits_opcode(wrapped_error_device_auto_buffer_in_d_bits_opcode),
    .auto_buffer_in_d_bits_size(wrapped_error_device_auto_buffer_in_d_bits_size),
    .auto_buffer_in_d_bits_source(wrapped_error_device_auto_buffer_in_d_bits_source),
    .auto_buffer_in_d_bits_denied(wrapped_error_device_auto_buffer_in_d_bits_denied),
    .auto_buffer_in_d_bits_data(wrapped_error_device_auto_buffer_in_d_bits_data),
    .auto_buffer_in_d_bits_corrupt(wrapped_error_device_auto_buffer_in_d_bits_corrupt),
    .io_covSum(wrapped_error_device_io_covSum)
  );
  TLInterconnectCoupler_7 coupler_to_plic ( // @[LazyModule.scala 432:27]
    .clock(coupler_to_plic_clock),
    .reset(coupler_to_plic_reset),
    .auto_fragmenter_out_a_ready(coupler_to_plic_auto_fragmenter_out_a_ready),
    .auto_fragmenter_out_a_valid(coupler_to_plic_auto_fragmenter_out_a_valid),
    .auto_fragmenter_out_a_bits_opcode(coupler_to_plic_auto_fragmenter_out_a_bits_opcode),
    .auto_fragmenter_out_a_bits_size(coupler_to_plic_auto_fragmenter_out_a_bits_size),
    .auto_fragmenter_out_a_bits_source(coupler_to_plic_auto_fragmenter_out_a_bits_source),
    .auto_fragmenter_out_a_bits_address(coupler_to_plic_auto_fragmenter_out_a_bits_address),
    .auto_fragmenter_out_a_bits_mask(coupler_to_plic_auto_fragmenter_out_a_bits_mask),
    .auto_fragmenter_out_a_bits_data(coupler_to_plic_auto_fragmenter_out_a_bits_data),
    .auto_fragmenter_out_d_ready(coupler_to_plic_auto_fragmenter_out_d_ready),
    .auto_fragmenter_out_d_valid(coupler_to_plic_auto_fragmenter_out_d_valid),
    .auto_fragmenter_out_d_bits_opcode(coupler_to_plic_auto_fragmenter_out_d_bits_opcode),
    .auto_fragmenter_out_d_bits_size(coupler_to_plic_auto_fragmenter_out_d_bits_size),
    .auto_fragmenter_out_d_bits_source(coupler_to_plic_auto_fragmenter_out_d_bits_source),
    .auto_fragmenter_out_d_bits_data(coupler_to_plic_auto_fragmenter_out_d_bits_data),
    .auto_tl_in_a_ready(coupler_to_plic_auto_tl_in_a_ready),
    .auto_tl_in_a_valid(coupler_to_plic_auto_tl_in_a_valid),
    .auto_tl_in_a_bits_opcode(coupler_to_plic_auto_tl_in_a_bits_opcode),
    .auto_tl_in_a_bits_size(coupler_to_plic_auto_tl_in_a_bits_size),
    .auto_tl_in_a_bits_source(coupler_to_plic_auto_tl_in_a_bits_source),
    .auto_tl_in_a_bits_address(coupler_to_plic_auto_tl_in_a_bits_address),
    .auto_tl_in_a_bits_mask(coupler_to_plic_auto_tl_in_a_bits_mask),
    .auto_tl_in_a_bits_data(coupler_to_plic_auto_tl_in_a_bits_data),
    .auto_tl_in_d_ready(coupler_to_plic_auto_tl_in_d_ready),
    .auto_tl_in_d_valid(coupler_to_plic_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_opcode(coupler_to_plic_auto_tl_in_d_bits_opcode),
    .auto_tl_in_d_bits_size(coupler_to_plic_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source(coupler_to_plic_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_data(coupler_to_plic_auto_tl_in_d_bits_data),
    .io_covSum(coupler_to_plic_io_covSum),
    .metaReset(coupler_to_plic_metaReset)
  );
  TLInterconnectCoupler_8 coupler_to_clint ( // @[LazyModule.scala 432:27]
    .clock(coupler_to_clint_clock),
    .reset(coupler_to_clint_reset),
    .auto_fragmenter_out_a_ready(coupler_to_clint_auto_fragmenter_out_a_ready),
    .auto_fragmenter_out_a_valid(coupler_to_clint_auto_fragmenter_out_a_valid),
    .auto_fragmenter_out_a_bits_opcode(coupler_to_clint_auto_fragmenter_out_a_bits_opcode),
    .auto_fragmenter_out_a_bits_size(coupler_to_clint_auto_fragmenter_out_a_bits_size),
    .auto_fragmenter_out_a_bits_source(coupler_to_clint_auto_fragmenter_out_a_bits_source),
    .auto_fragmenter_out_a_bits_address(coupler_to_clint_auto_fragmenter_out_a_bits_address),
    .auto_fragmenter_out_a_bits_mask(coupler_to_clint_auto_fragmenter_out_a_bits_mask),
    .auto_fragmenter_out_a_bits_data(coupler_to_clint_auto_fragmenter_out_a_bits_data),
    .auto_fragmenter_out_d_ready(coupler_to_clint_auto_fragmenter_out_d_ready),
    .auto_fragmenter_out_d_valid(coupler_to_clint_auto_fragmenter_out_d_valid),
    .auto_fragmenter_out_d_bits_opcode(coupler_to_clint_auto_fragmenter_out_d_bits_opcode),
    .auto_fragmenter_out_d_bits_size(coupler_to_clint_auto_fragmenter_out_d_bits_size),
    .auto_fragmenter_out_d_bits_source(coupler_to_clint_auto_fragmenter_out_d_bits_source),
    .auto_fragmenter_out_d_bits_data(coupler_to_clint_auto_fragmenter_out_d_bits_data),
    .auto_tl_in_a_ready(coupler_to_clint_auto_tl_in_a_ready),
    .auto_tl_in_a_valid(coupler_to_clint_auto_tl_in_a_valid),
    .auto_tl_in_a_bits_opcode(coupler_to_clint_auto_tl_in_a_bits_opcode),
    .auto_tl_in_a_bits_size(coupler_to_clint_auto_tl_in_a_bits_size),
    .auto_tl_in_a_bits_source(coupler_to_clint_auto_tl_in_a_bits_source),
    .auto_tl_in_a_bits_address(coupler_to_clint_auto_tl_in_a_bits_address),
    .auto_tl_in_a_bits_mask(coupler_to_clint_auto_tl_in_a_bits_mask),
    .auto_tl_in_a_bits_data(coupler_to_clint_auto_tl_in_a_bits_data),
    .auto_tl_in_d_ready(coupler_to_clint_auto_tl_in_d_ready),
    .auto_tl_in_d_valid(coupler_to_clint_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_opcode(coupler_to_clint_auto_tl_in_d_bits_opcode),
    .auto_tl_in_d_bits_size(coupler_to_clint_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source(coupler_to_clint_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_data(coupler_to_clint_auto_tl_in_d_bits_data),
    .io_covSum(coupler_to_clint_io_covSum),
    .metaReset(coupler_to_clint_metaReset)
  );
  TLInterconnectCoupler_10 coupler_to_bootrom ( // @[LazyModule.scala 432:27]
    .clock(coupler_to_bootrom_clock),
    .reset(coupler_to_bootrom_reset),
    .auto_fragmenter_out_a_ready(coupler_to_bootrom_auto_fragmenter_out_a_ready),
    .auto_fragmenter_out_a_valid(coupler_to_bootrom_auto_fragmenter_out_a_valid),
    .auto_fragmenter_out_a_bits_size(coupler_to_bootrom_auto_fragmenter_out_a_bits_size),
    .auto_fragmenter_out_a_bits_source(coupler_to_bootrom_auto_fragmenter_out_a_bits_source),
    .auto_fragmenter_out_a_bits_address(coupler_to_bootrom_auto_fragmenter_out_a_bits_address),
    .auto_fragmenter_out_d_ready(coupler_to_bootrom_auto_fragmenter_out_d_ready),
    .auto_fragmenter_out_d_valid(coupler_to_bootrom_auto_fragmenter_out_d_valid),
    .auto_fragmenter_out_d_bits_size(coupler_to_bootrom_auto_fragmenter_out_d_bits_size),
    .auto_fragmenter_out_d_bits_source(coupler_to_bootrom_auto_fragmenter_out_d_bits_source),
    .auto_fragmenter_out_d_bits_data(coupler_to_bootrom_auto_fragmenter_out_d_bits_data),
    .auto_tl_in_a_ready(coupler_to_bootrom_auto_tl_in_a_ready),
    .auto_tl_in_a_valid(coupler_to_bootrom_auto_tl_in_a_valid),
    .auto_tl_in_a_bits_size(coupler_to_bootrom_auto_tl_in_a_bits_size),
    .auto_tl_in_a_bits_source(coupler_to_bootrom_auto_tl_in_a_bits_source),
    .auto_tl_in_a_bits_address(coupler_to_bootrom_auto_tl_in_a_bits_address),
    .auto_tl_in_a_bits_mask(coupler_to_bootrom_auto_tl_in_a_bits_mask),
    .auto_tl_in_d_ready(coupler_to_bootrom_auto_tl_in_d_ready),
    .auto_tl_in_d_valid(coupler_to_bootrom_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_size(coupler_to_bootrom_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source(coupler_to_bootrom_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_data(coupler_to_bootrom_auto_tl_in_d_bits_data),
    .io_covSum(coupler_to_bootrom_io_covSum),
    .metaReset(coupler_to_bootrom_metaReset)
  );
  TLInterconnectCoupler_11 coupler_to_MaskROM ( // @[LazyModule.scala 432:27]
    .clock(coupler_to_MaskROM_clock),
    .reset(coupler_to_MaskROM_reset),
    .auto_fragmenter_out_a_ready(coupler_to_MaskROM_auto_fragmenter_out_a_ready),
    .auto_fragmenter_out_a_valid(coupler_to_MaskROM_auto_fragmenter_out_a_valid),
    .auto_fragmenter_out_a_bits_size(coupler_to_MaskROM_auto_fragmenter_out_a_bits_size),
    .auto_fragmenter_out_a_bits_source(coupler_to_MaskROM_auto_fragmenter_out_a_bits_source),
    .auto_fragmenter_out_a_bits_address(coupler_to_MaskROM_auto_fragmenter_out_a_bits_address),
    .auto_fragmenter_out_d_ready(coupler_to_MaskROM_auto_fragmenter_out_d_ready),
    .auto_fragmenter_out_d_valid(coupler_to_MaskROM_auto_fragmenter_out_d_valid),
    .auto_fragmenter_out_d_bits_size(coupler_to_MaskROM_auto_fragmenter_out_d_bits_size),
    .auto_fragmenter_out_d_bits_source(coupler_to_MaskROM_auto_fragmenter_out_d_bits_source),
    .auto_fragmenter_out_d_bits_data(coupler_to_MaskROM_auto_fragmenter_out_d_bits_data),
    .auto_tl_in_a_ready(coupler_to_MaskROM_auto_tl_in_a_ready),
    .auto_tl_in_a_valid(coupler_to_MaskROM_auto_tl_in_a_valid),
    .auto_tl_in_a_bits_size(coupler_to_MaskROM_auto_tl_in_a_bits_size),
    .auto_tl_in_a_bits_source(coupler_to_MaskROM_auto_tl_in_a_bits_source),
    .auto_tl_in_a_bits_address(coupler_to_MaskROM_auto_tl_in_a_bits_address),
    .auto_tl_in_a_bits_mask(coupler_to_MaskROM_auto_tl_in_a_bits_mask),
    .auto_tl_in_d_ready(coupler_to_MaskROM_auto_tl_in_d_ready),
    .auto_tl_in_d_valid(coupler_to_MaskROM_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_size(coupler_to_MaskROM_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source(coupler_to_MaskROM_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_data(coupler_to_MaskROM_auto_tl_in_d_bits_data),
    .io_covSum(coupler_to_MaskROM_io_covSum),
    .metaReset(coupler_to_MaskROM_metaReset)
  );
  TLInterconnectCoupler_12 coupler_to_magic ( // @[LazyModule.scala 432:27]
    .clock(coupler_to_magic_clock),
    .reset(coupler_to_magic_reset),
    .auto_fragmenter_out_a_ready(coupler_to_magic_auto_fragmenter_out_a_ready),
    .auto_fragmenter_out_a_valid(coupler_to_magic_auto_fragmenter_out_a_valid),
    .auto_fragmenter_out_a_bits_opcode(coupler_to_magic_auto_fragmenter_out_a_bits_opcode),
    .auto_fragmenter_out_a_bits_size(coupler_to_magic_auto_fragmenter_out_a_bits_size),
    .auto_fragmenter_out_a_bits_source(coupler_to_magic_auto_fragmenter_out_a_bits_source),
    .auto_fragmenter_out_a_bits_address(coupler_to_magic_auto_fragmenter_out_a_bits_address),
    .auto_fragmenter_out_a_bits_mask(coupler_to_magic_auto_fragmenter_out_a_bits_mask),
    .auto_fragmenter_out_d_ready(coupler_to_magic_auto_fragmenter_out_d_ready),
    .auto_fragmenter_out_d_valid(coupler_to_magic_auto_fragmenter_out_d_valid),
    .auto_fragmenter_out_d_bits_opcode(coupler_to_magic_auto_fragmenter_out_d_bits_opcode),
    .auto_fragmenter_out_d_bits_size(coupler_to_magic_auto_fragmenter_out_d_bits_size),
    .auto_fragmenter_out_d_bits_source(coupler_to_magic_auto_fragmenter_out_d_bits_source),
    .auto_fragmenter_out_d_bits_data(coupler_to_magic_auto_fragmenter_out_d_bits_data),
    .auto_tl_in_a_ready(coupler_to_magic_auto_tl_in_a_ready),
    .auto_tl_in_a_valid(coupler_to_magic_auto_tl_in_a_valid),
    .auto_tl_in_a_bits_opcode(coupler_to_magic_auto_tl_in_a_bits_opcode),
    .auto_tl_in_a_bits_size(coupler_to_magic_auto_tl_in_a_bits_size),
    .auto_tl_in_a_bits_source(coupler_to_magic_auto_tl_in_a_bits_source),
    .auto_tl_in_a_bits_address(coupler_to_magic_auto_tl_in_a_bits_address),
    .auto_tl_in_a_bits_mask(coupler_to_magic_auto_tl_in_a_bits_mask),
    .auto_tl_in_d_ready(coupler_to_magic_auto_tl_in_d_ready),
    .auto_tl_in_d_valid(coupler_to_magic_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_opcode(coupler_to_magic_auto_tl_in_d_bits_opcode),
    .auto_tl_in_d_bits_size(coupler_to_magic_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source(coupler_to_magic_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_data(coupler_to_magic_auto_tl_in_d_bits_data),
    .io_covSum(coupler_to_magic_io_covSum),
    .metaReset(coupler_to_magic_metaReset)
  );
  assign subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_clock =
    subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_reset =
    subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_clock =
    subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_reset =
    subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_clock = clockGroup_auto_in_member_subsystem_cbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_reset = clockGroup_auto_in_member_subsystem_cbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_in_a_ready = in_xbar_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_valid = in_xbar_auto_out_d_valid; // @[ReadyValidCancel.scala 21:38]
  assign in_xbar_auto_in_d_bits_opcode = in_xbar_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_bits_size = in_xbar_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_bits_source = in_xbar_auto_out_d_bits_source; // @[Xbar.scala 228:69]
  assign in_xbar_auto_in_d_bits_denied = in_xbar_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_bits_data = in_xbar_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_in_d_bits_corrupt = in_xbar_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign in_xbar_auto_out_a_valid = in_xbar_auto_in_a_valid; // @[ReadyValidCancel.scala 21:38]
  assign in_xbar_auto_out_a_bits_opcode = in_xbar_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_param = in_xbar_auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_size = in_xbar_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_source = in_xbar_auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign in_xbar_auto_out_a_bits_address = in_xbar_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_mask = in_xbar_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_a_bits_data = in_xbar_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_xbar_auto_out_d_ready = in_xbar_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_ready = buffer_1_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_in_d_valid = buffer_1_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_in_d_bits_opcode = buffer_1_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_in_d_bits_size = buffer_1_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_in_d_bits_source = buffer_1_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_in_d_bits_denied = buffer_1_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_in_d_bits_data = buffer_1_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_in_d_bits_corrupt = buffer_1_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_out_a_valid = buffer_1_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_a_bits_opcode = buffer_1_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_a_bits_param = buffer_1_auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_a_bits_size = buffer_1_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_a_bits_source = buffer_1_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_a_bits_address = buffer_1_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_a_bits_mask = buffer_1_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_a_bits_data = buffer_1_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_d_ready = buffer_1_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_ready =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_valid =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_opcode =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_size =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_source =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_denied =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_data =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_corrupt =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_valid =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_param =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_size =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_source =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_address =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_mask =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_data =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_ready =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_ready =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_ready; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_valid =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_valid; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_opcode =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_size =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_source =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_denied =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_denied; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_data =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_corrupt =
    coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_valid =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_param =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_size =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_source =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_address =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_mask =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_data =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_ready =
    coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_valid =
    coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_valid; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_opcode =
    coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_param =
    coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_param; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_size =
    coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_source =
    coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_address =
    coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_mask =
    coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_a_bits_data =
    coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_in_d_ready =
    coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_ready; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_a_ready =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_valid =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_opcode =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_size =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_source =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_denied =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_data =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_widget_auto_out_d_bits_corrupt =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_coupler_to_magic_fragmenter_out_a_valid = coupler_to_magic_auto_fragmenter_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_magic_fragmenter_out_a_bits_opcode = coupler_to_magic_auto_fragmenter_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_magic_fragmenter_out_a_bits_size = coupler_to_magic_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_magic_fragmenter_out_a_bits_source = coupler_to_magic_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_magic_fragmenter_out_a_bits_address = coupler_to_magic_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_magic_fragmenter_out_a_bits_mask = coupler_to_magic_auto_fragmenter_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_magic_fragmenter_out_d_ready = coupler_to_magic_auto_fragmenter_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_MaskROM_fragmenter_out_a_valid = coupler_to_MaskROM_auto_fragmenter_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_MaskROM_fragmenter_out_a_bits_size = coupler_to_MaskROM_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_MaskROM_fragmenter_out_a_bits_source = coupler_to_MaskROM_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_MaskROM_fragmenter_out_a_bits_address = coupler_to_MaskROM_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_MaskROM_fragmenter_out_d_ready = coupler_to_MaskROM_auto_fragmenter_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bootrom_fragmenter_out_a_valid = coupler_to_bootrom_auto_fragmenter_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bootrom_fragmenter_out_a_bits_size = coupler_to_bootrom_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bootrom_fragmenter_out_a_bits_source = coupler_to_bootrom_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bootrom_fragmenter_out_a_bits_address = coupler_to_bootrom_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bootrom_fragmenter_out_d_ready = coupler_to_bootrom_auto_fragmenter_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_clint_fragmenter_out_a_valid = coupler_to_clint_auto_fragmenter_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_clint_fragmenter_out_a_bits_opcode = coupler_to_clint_auto_fragmenter_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_clint_fragmenter_out_a_bits_size = coupler_to_clint_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_clint_fragmenter_out_a_bits_source = coupler_to_clint_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_clint_fragmenter_out_a_bits_address = coupler_to_clint_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_clint_fragmenter_out_a_bits_mask = coupler_to_clint_auto_fragmenter_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_clint_fragmenter_out_a_bits_data = coupler_to_clint_auto_fragmenter_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_clint_fragmenter_out_d_ready = coupler_to_clint_auto_fragmenter_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_plic_fragmenter_out_a_valid = coupler_to_plic_auto_fragmenter_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_plic_fragmenter_out_a_bits_opcode = coupler_to_plic_auto_fragmenter_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_plic_fragmenter_out_a_bits_size = coupler_to_plic_auto_fragmenter_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_plic_fragmenter_out_a_bits_source = coupler_to_plic_auto_fragmenter_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_plic_fragmenter_out_a_bits_address = coupler_to_plic_auto_fragmenter_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_plic_fragmenter_out_a_bits_mask = coupler_to_plic_auto_fragmenter_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_plic_fragmenter_out_a_bits_data = coupler_to_plic_auto_fragmenter_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_plic_fragmenter_out_d_ready = coupler_to_plic_auto_fragmenter_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_param; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready =
    coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_fixedClockNode_out_0_clock = fixedClockNode_auto_out_1_clock; // @[LazyModule.scala 311:12]
  assign auto_fixedClockNode_out_0_reset = fixedClockNode_auto_out_1_reset; // @[LazyModule.scala 311:12]
  assign auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock =
    subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_clock; // @[LazyModule.scala 311:12]
  assign auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset =
    subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_reset; // @[LazyModule.scala 311:12]
  assign auto_bus_xing_in_a_ready = buffer_1_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_valid = buffer_1_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_opcode = buffer_1_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_size = buffer_1_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_source = buffer_1_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_denied = buffer_1_auto_in_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_data = buffer_1_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_corrupt = buffer_1_auto_in_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_clock =
    auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock; // @[LazyModule.scala 309:16]
  assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_reset =
    auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset; // @[LazyModule.scala 309:16]
  assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_clock =
    auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock; // @[LazyModule.scala 309:16]
  assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_reset =
    auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset; // @[LazyModule.scala 309:16]
  assign clockGroup_auto_in_member_subsystem_cbus_0_clock =
    subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_clock; // @[LazyModule.scala 298:16]
  assign clockGroup_auto_in_member_subsystem_cbus_0_reset =
    subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_reset; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[LazyModule.scala 298:16]
  assign fixer_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign fixer_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign fixer_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_param = buffer_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_a_ready = out_xbar_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_valid = out_xbar_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_opcode = out_xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_size = out_xbar_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_source = out_xbar_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_denied = out_xbar_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_data = out_xbar_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign fixer_auto_out_d_bits_corrupt = out_xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_in_a_valid = buffer_1_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_param = buffer_1_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_size = buffer_1_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_source = buffer_1_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_address = buffer_1_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_mask = buffer_1_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_a_bits_data = buffer_1_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_in_d_ready = buffer_1_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign in_xbar_auto_out_a_ready = atomics_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_valid = atomics_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_opcode = atomics_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_size = atomics_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_source = atomics_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_denied = atomics_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_data = atomics_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign in_xbar_auto_out_d_bits_corrupt = atomics_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign out_xbar_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign out_xbar_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign out_xbar_auto_in_a_valid = fixer_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_param = fixer_auto_out_a_bits_param; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_size = fixer_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_source = fixer_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_address = fixer_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_a_bits_data = fixer_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_in_d_ready = fixer_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_6_a_ready = coupler_to_magic_auto_tl_in_a_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_6_d_valid = coupler_to_magic_auto_tl_in_d_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_6_d_bits_opcode = coupler_to_magic_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_6_d_bits_size = coupler_to_magic_auto_tl_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_6_d_bits_source = coupler_to_magic_auto_tl_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_6_d_bits_data = coupler_to_magic_auto_tl_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_5_a_ready = coupler_to_MaskROM_auto_tl_in_a_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_5_d_valid = coupler_to_MaskROM_auto_tl_in_d_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_5_d_bits_size = coupler_to_MaskROM_auto_tl_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_5_d_bits_source = coupler_to_MaskROM_auto_tl_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_5_d_bits_data = coupler_to_MaskROM_auto_tl_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_4_a_ready = coupler_to_bootrom_auto_tl_in_a_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_4_d_valid = coupler_to_bootrom_auto_tl_in_d_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_4_d_bits_size = coupler_to_bootrom_auto_tl_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_4_d_bits_source = coupler_to_bootrom_auto_tl_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_4_d_bits_data = coupler_to_bootrom_auto_tl_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_3_a_ready = coupler_to_clint_auto_tl_in_a_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_3_d_valid = coupler_to_clint_auto_tl_in_d_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_3_d_bits_opcode = coupler_to_clint_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_3_d_bits_size = coupler_to_clint_auto_tl_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_3_d_bits_source = coupler_to_clint_auto_tl_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_3_d_bits_data = coupler_to_clint_auto_tl_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_2_a_ready = coupler_to_plic_auto_tl_in_a_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_2_d_valid = coupler_to_plic_auto_tl_in_d_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_2_d_bits_opcode = coupler_to_plic_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_2_d_bits_size = coupler_to_plic_auto_tl_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_2_d_bits_source = coupler_to_plic_auto_tl_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_2_d_bits_data = coupler_to_plic_auto_tl_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_1_a_ready = coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_1_d_valid = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_1_d_bits_opcode = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_1_d_bits_size = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_1_d_bits_source = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_1_d_bits_denied = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_1_d_bits_data = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_1_d_bits_corrupt = coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_0_a_ready = wrapped_error_device_auto_buffer_in_a_ready; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_0_d_valid = wrapped_error_device_auto_buffer_in_d_valid; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_0_d_bits_opcode = wrapped_error_device_auto_buffer_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_0_d_bits_size = wrapped_error_device_auto_buffer_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_0_d_bits_source = wrapped_error_device_auto_buffer_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_0_d_bits_denied = wrapped_error_device_auto_buffer_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_0_d_bits_data = wrapped_error_device_auto_buffer_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign out_xbar_auto_out_0_d_bits_corrupt = wrapped_error_device_auto_buffer_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign buffer_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign buffer_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign buffer_auto_in_a_valid = atomics_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_opcode = atomics_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_param = atomics_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_size = atomics_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_source = atomics_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_address = atomics_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_mask = atomics_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_data = atomics_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_d_ready = atomics_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_a_ready = fixer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_valid = fixer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_size = fixer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_source = fixer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_denied = fixer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_data = fixer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign atomics_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign atomics_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign atomics_auto_in_a_valid = in_xbar_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_opcode = in_xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_param = in_xbar_auto_out_a_bits_param; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_size = in_xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_source = in_xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_address = in_xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_mask = in_xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_a_bits_data = in_xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign atomics_auto_in_d_ready = in_xbar_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign atomics_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign atomics_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign wrapped_error_device_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign wrapped_error_device_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign wrapped_error_device_auto_buffer_in_a_valid = out_xbar_auto_out_0_a_valid; // @[LazyModule.scala 298:16]
  assign wrapped_error_device_auto_buffer_in_a_bits_opcode = out_xbar_auto_out_0_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign wrapped_error_device_auto_buffer_in_a_bits_size = out_xbar_auto_out_0_a_bits_size; // @[LazyModule.scala 298:16]
  assign wrapped_error_device_auto_buffer_in_a_bits_source = out_xbar_auto_out_0_a_bits_source; // @[LazyModule.scala 298:16]
  assign wrapped_error_device_auto_buffer_in_d_ready = out_xbar_auto_out_0_d_ready; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_valid = auto_bus_xing_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_opcode = auto_bus_xing_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_param = auto_bus_xing_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_size = auto_bus_xing_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_source = auto_bus_xing_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_address = auto_bus_xing_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_mask = auto_bus_xing_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_bits_data = auto_bus_xing_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_d_ready = auto_bus_xing_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_out_a_ready = in_xbar_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_valid = in_xbar_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_opcode = in_xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_size = in_xbar_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_source = in_xbar_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_denied = in_xbar_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_data = in_xbar_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign buffer_1_auto_out_d_bits_corrupt = in_xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_valid = out_xbar_auto_out_1_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_opcode = out_xbar_auto_out_1_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_param = out_xbar_auto_out_1_a_bits_param; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_size = out_xbar_auto_out_1_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_source = out_xbar_auto_out_1_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_address = out_xbar_auto_out_1_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_mask = out_xbar_auto_out_1_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_a_bits_data = out_xbar_auto_out_1_a_bits_data; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_widget_in_d_ready = out_xbar_auto_out_1_d_ready; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_a_ready =
    auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_valid =
    auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_opcode =
    auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_size =
    auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_source =
    auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_denied =
    auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_data =
    auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_pbus_auto_bus_xing_out_d_bits_corrupt =
    auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign coupler_to_plic_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_plic_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_plic_auto_fragmenter_out_a_ready = auto_coupler_to_plic_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_plic_auto_fragmenter_out_d_valid = auto_coupler_to_plic_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_plic_auto_fragmenter_out_d_bits_opcode = auto_coupler_to_plic_fragmenter_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_plic_auto_fragmenter_out_d_bits_size = auto_coupler_to_plic_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_plic_auto_fragmenter_out_d_bits_source = auto_coupler_to_plic_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_plic_auto_fragmenter_out_d_bits_data = auto_coupler_to_plic_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_plic_auto_tl_in_a_valid = out_xbar_auto_out_2_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_plic_auto_tl_in_a_bits_opcode = out_xbar_auto_out_2_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign coupler_to_plic_auto_tl_in_a_bits_size = out_xbar_auto_out_2_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_plic_auto_tl_in_a_bits_source = out_xbar_auto_out_2_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_plic_auto_tl_in_a_bits_address = out_xbar_auto_out_2_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_plic_auto_tl_in_a_bits_mask = out_xbar_auto_out_2_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_plic_auto_tl_in_a_bits_data = out_xbar_auto_out_2_a_bits_data; // @[LazyModule.scala 298:16]
  assign coupler_to_plic_auto_tl_in_d_ready = out_xbar_auto_out_2_d_ready; // @[LazyModule.scala 298:16]
  assign coupler_to_clint_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_clint_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_clint_auto_fragmenter_out_a_ready = auto_coupler_to_clint_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_clint_auto_fragmenter_out_d_valid = auto_coupler_to_clint_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_clint_auto_fragmenter_out_d_bits_opcode = auto_coupler_to_clint_fragmenter_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_clint_auto_fragmenter_out_d_bits_size = auto_coupler_to_clint_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_clint_auto_fragmenter_out_d_bits_source = auto_coupler_to_clint_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_clint_auto_fragmenter_out_d_bits_data = auto_coupler_to_clint_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_clint_auto_tl_in_a_valid = out_xbar_auto_out_3_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_clint_auto_tl_in_a_bits_opcode = out_xbar_auto_out_3_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign coupler_to_clint_auto_tl_in_a_bits_size = out_xbar_auto_out_3_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_clint_auto_tl_in_a_bits_source = out_xbar_auto_out_3_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_clint_auto_tl_in_a_bits_address = out_xbar_auto_out_3_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_clint_auto_tl_in_a_bits_mask = out_xbar_auto_out_3_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_clint_auto_tl_in_a_bits_data = out_xbar_auto_out_3_a_bits_data; // @[LazyModule.scala 298:16]
  assign coupler_to_clint_auto_tl_in_d_ready = out_xbar_auto_out_3_d_ready; // @[LazyModule.scala 298:16]
  assign coupler_to_bootrom_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bootrom_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bootrom_auto_fragmenter_out_a_ready = auto_coupler_to_bootrom_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_bootrom_auto_fragmenter_out_d_valid = auto_coupler_to_bootrom_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_bootrom_auto_fragmenter_out_d_bits_size = auto_coupler_to_bootrom_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_bootrom_auto_fragmenter_out_d_bits_source = auto_coupler_to_bootrom_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_bootrom_auto_fragmenter_out_d_bits_data = auto_coupler_to_bootrom_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_bootrom_auto_tl_in_a_valid = out_xbar_auto_out_4_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_bootrom_auto_tl_in_a_bits_size = out_xbar_auto_out_4_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_bootrom_auto_tl_in_a_bits_source = out_xbar_auto_out_4_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_bootrom_auto_tl_in_a_bits_address = out_xbar_auto_out_4_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_bootrom_auto_tl_in_a_bits_mask = out_xbar_auto_out_4_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_bootrom_auto_tl_in_d_ready = out_xbar_auto_out_4_d_ready; // @[LazyModule.scala 298:16]
  assign coupler_to_MaskROM_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_MaskROM_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_MaskROM_auto_fragmenter_out_a_ready = auto_coupler_to_MaskROM_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_MaskROM_auto_fragmenter_out_d_valid = auto_coupler_to_MaskROM_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_MaskROM_auto_fragmenter_out_d_bits_size = auto_coupler_to_MaskROM_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_MaskROM_auto_fragmenter_out_d_bits_source = auto_coupler_to_MaskROM_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_MaskROM_auto_fragmenter_out_d_bits_data = auto_coupler_to_MaskROM_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_MaskROM_auto_tl_in_a_valid = out_xbar_auto_out_5_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_MaskROM_auto_tl_in_a_bits_size = out_xbar_auto_out_5_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_MaskROM_auto_tl_in_a_bits_source = out_xbar_auto_out_5_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_MaskROM_auto_tl_in_a_bits_address = out_xbar_auto_out_5_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_MaskROM_auto_tl_in_a_bits_mask = out_xbar_auto_out_5_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_MaskROM_auto_tl_in_d_ready = out_xbar_auto_out_5_d_ready; // @[LazyModule.scala 298:16]
  assign coupler_to_magic_clock = fixedClockNode_auto_out_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_magic_reset = fixedClockNode_auto_out_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_magic_auto_fragmenter_out_a_ready = auto_coupler_to_magic_fragmenter_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_magic_auto_fragmenter_out_d_valid = auto_coupler_to_magic_fragmenter_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_magic_auto_fragmenter_out_d_bits_opcode = auto_coupler_to_magic_fragmenter_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_magic_auto_fragmenter_out_d_bits_size = auto_coupler_to_magic_fragmenter_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_magic_auto_fragmenter_out_d_bits_source = auto_coupler_to_magic_fragmenter_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_magic_auto_fragmenter_out_d_bits_data = auto_coupler_to_magic_fragmenter_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_magic_auto_tl_in_a_valid = out_xbar_auto_out_6_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_magic_auto_tl_in_a_bits_opcode = out_xbar_auto_out_6_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign coupler_to_magic_auto_tl_in_a_bits_size = out_xbar_auto_out_6_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_magic_auto_tl_in_a_bits_source = out_xbar_auto_out_6_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_magic_auto_tl_in_a_bits_address = out_xbar_auto_out_6_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_magic_auto_tl_in_a_bits_mask = out_xbar_auto_out_6_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_magic_auto_tl_in_d_ready = out_xbar_auto_out_6_d_ready; // @[LazyModule.scala 298:16]
  assign PeripheryBus_1_covSum = 30'h0;
  assign atomics_sum = PeripheryBus_1_covSum + atomics_io_covSum;
  assign coupler_to_clint_sum = atomics_sum + coupler_to_clint_io_covSum;
  assign wrapped_error_device_sum = coupler_to_clint_sum + wrapped_error_device_io_covSum;
  assign fixedClockNode_sum = wrapped_error_device_sum + fixedClockNode_io_covSum;
  assign fixer_sum = fixedClockNode_sum + fixer_io_covSum;
  assign coupler_to_bootrom_sum = fixer_sum + coupler_to_bootrom_io_covSum;
  assign out_xbar_sum = coupler_to_bootrom_sum + out_xbar_io_covSum;
  assign coupler_to_magic_sum = out_xbar_sum + coupler_to_magic_io_covSum;
  assign coupler_to_plic_sum = coupler_to_magic_sum + coupler_to_plic_io_covSum;
  assign coupler_to_MaskROM_sum = coupler_to_plic_sum + coupler_to_MaskROM_io_covSum;
  assign buffer_sum = coupler_to_MaskROM_sum + buffer_io_covSum;
  assign io_covSum = buffer_sum;
  assign atomics_metaReset = metaReset;
  assign coupler_to_clint_metaReset = metaReset;
  assign fixer_metaReset = metaReset;
  assign coupler_to_bootrom_metaReset = metaReset;
  assign out_xbar_metaReset = metaReset;
  assign coupler_to_magic_metaReset = metaReset;
  assign coupler_to_plic_metaReset = metaReset;
  assign coupler_to_MaskROM_metaReset = metaReset;
endmodule
module TLFIFOFixer_4(
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [8:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input         auto_in_a_bits_user_amba_prot_bufferable,
  input         auto_in_a_bits_user_amba_prot_modifiable,
  input         auto_in_a_bits_user_amba_prot_readalloc,
  input         auto_in_a_bits_user_amba_prot_writealloc,
  input         auto_in_a_bits_user_amba_prot_privileged,
  input         auto_in_a_bits_user_amba_prot_secure,
  input         auto_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [8:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_size,
  output [8:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output        auto_out_a_bits_user_amba_prot_bufferable,
  output        auto_out_a_bits_user_amba_prot_modifiable,
  output        auto_out_a_bits_user_amba_prot_readalloc,
  output        auto_out_a_bits_user_amba_prot_writealloc,
  output        auto_out_a_bits_user_amba_prot_privileged,
  output        auto_out_a_bits_user_amba_prot_secure,
  output        auto_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [2:0]  auto_out_d_bits_size,
  input  [8:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum
);
  wire [29:0] TLFIFOFixer_4_covSum;
  assign auto_in_a_ready = auto_out_a_ready; // @[FIFOFixer.scala 88:33]
  assign auto_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[FIFOFixer.scala 87:33]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLFIFOFixer_4_covSum = 30'h0;
  assign io_covSum = TLFIFOFixer_4_covSum;
endmodule
module ProbePicker(
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [8:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input         auto_in_a_bits_user_amba_prot_bufferable,
  input         auto_in_a_bits_user_amba_prot_modifiable,
  input         auto_in_a_bits_user_amba_prot_readalloc,
  input         auto_in_a_bits_user_amba_prot_writealloc,
  input         auto_in_a_bits_user_amba_prot_privileged,
  input         auto_in_a_bits_user_amba_prot_secure,
  input         auto_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [8:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_size,
  output [8:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output        auto_out_a_bits_user_amba_prot_bufferable,
  output        auto_out_a_bits_user_amba_prot_modifiable,
  output        auto_out_a_bits_user_amba_prot_readalloc,
  output        auto_out_a_bits_user_amba_prot_writealloc,
  output        auto_out_a_bits_user_amba_prot_privileged,
  output        auto_out_a_bits_user_amba_prot_secure,
  output        auto_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [2:0]  auto_out_d_bits_size,
  input  [8:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum
);
  wire [29:0] ProbePicker_covSum;
  assign auto_in_a_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign ProbePicker_covSum = 30'h0;
  assign io_covSum = ProbePicker_covSum;
endmodule
module QueueCompatibility_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_tl_state_size,
  input  [8:0]  io_enq_bits_tl_state_source,
  input  [4:0]  io_enq_bits_extra_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_tl_state_size,
  output [8:0]  io_deq_bits_tl_state_source,
  output [4:0]  io_deq_bits_extra_id,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:31]; // @[Decoupled.scala 259:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [4:0] ram_tl_state_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_tl_state_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_tl_state_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_tl_state_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [8:0] ram_tl_state_source [0:31]; // @[Decoupled.scala 259:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [4:0] ram_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [8:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [8:0] ram_tl_state_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_tl_state_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_tl_state_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_tl_state_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] ram_extra_id [0:31]; // @[Decoupled.scala 259:95]
  wire  ram_extra_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [4:0] ram_extra_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [4:0] ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_extra_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_extra_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_extra_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_extra_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [4:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [4:0] _value_T_1 = enq_ptr_value + 5'h1; // @[Counter.scala 78:24]
  wire [4:0] _value_T_3 = deq_ptr_value + 5'h1; // @[Counter.scala 78:24]
  wire [29:0] QueueCompatibility_4_covSum;
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = enq_ptr_value;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = enq_ptr_value;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_extra_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_extra_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_extra_id_io_deq_bits_MPORT_data = ram_extra_id[ram_extra_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_extra_id_MPORT_data = io_enq_bits_extra_id;
  assign ram_extra_id_MPORT_addr = enq_ptr_value;
  assign ram_extra_id_MPORT_mask = 1'h1;
  assign ram_extra_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_extra_id = ram_extra_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign QueueCompatibility_4_covSum = 30'h0;
  assign io_covSum = QueueCompatibility_4_covSum;
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_extra_id_MPORT_en & ram_extra_id_MPORT_mask) begin
      ram_extra_id[ram_extra_id_MPORT_addr] <= ram_extra_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 5'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      enq_ptr_value <= _value_T_1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 5'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      deq_ptr_value <= _value_T_3;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram_extra_id[initvar] = _RAND_2[4:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4UserYanker_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  input  [3:0]  auto_in_aw_bits_echo_tl_state_size,
  input  [8:0]  auto_in_aw_bits_echo_tl_state_source,
  input  [4:0]  auto_in_aw_bits_echo_extra_id,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [3:0]  auto_in_b_bits_echo_tl_state_size,
  output [8:0]  auto_in_b_bits_echo_tl_state_source,
  output [4:0]  auto_in_b_bits_echo_extra_id,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input  [3:0]  auto_in_ar_bits_echo_tl_state_size,
  input  [8:0]  auto_in_ar_bits_echo_tl_state_source,
  input  [4:0]  auto_in_ar_bits_echo_extra_id,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [3:0]  auto_in_r_bits_echo_tl_state_size,
  output [8:0]  auto_in_r_bits_echo_tl_state_source,
  output [4:0]  auto_in_r_bits_echo_extra_id,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last,
  output [29:0] io_covSum
);
  wire  QueueCompatibility_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_1_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_1_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_1_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_1_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_1_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_1_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_2_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_2_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_2_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_2_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_2_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_2_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_3_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_3_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_3_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_3_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_3_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_3_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_4_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_4_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_4_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_4_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_4_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_4_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_5_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_5_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_5_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_5_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_5_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_5_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_6_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_6_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_6_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_6_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_6_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_6_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_7_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_7_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_7_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_7_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_7_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_7_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_8_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_8_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_8_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_8_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_8_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_8_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_8_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_9_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_9_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_9_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_9_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_9_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_9_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_9_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_10_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_10_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_10_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_10_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_10_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_10_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_10_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_11_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_11_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_11_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_11_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_11_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_11_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_11_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_12_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_12_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_12_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_12_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_12_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_12_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_12_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_13_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_13_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_13_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_13_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_13_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_13_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_13_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_14_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_14_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_14_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_14_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_14_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_14_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_14_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_15_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_15_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_15_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_15_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_15_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_15_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_15_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_16_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_16_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_16_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_16_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_16_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_16_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_16_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_17_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_17_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_17_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_17_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_17_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_17_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_17_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_18_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_18_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_18_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_18_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_18_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_18_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_18_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_19_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_19_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_19_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_19_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_19_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_19_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_19_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_20_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_20_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_20_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_20_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_20_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_20_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_20_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_21_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_21_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_21_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_21_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_21_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_21_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_21_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_22_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_22_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_22_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_22_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_22_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_22_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_22_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_23_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_23_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_23_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_23_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_23_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_23_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_23_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_24_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_24_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_24_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_24_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_24_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_24_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_24_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_25_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_25_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_25_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_25_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_25_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_25_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_25_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_26_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_26_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_26_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_26_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_26_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_26_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_26_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_27_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_27_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_27_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_27_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_27_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_27_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_27_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_28_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_28_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_28_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_28_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_28_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_28_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_28_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_29_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_29_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_29_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_29_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_29_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_29_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_29_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_30_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_30_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_30_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_30_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_30_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_30_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_30_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_enq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_31_io_enq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_31_io_enq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_31_io_enq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_deq_valid; // @[UserYanker.scala 47:17]
  wire [3:0] QueueCompatibility_31_io_deq_bits_tl_state_size; // @[UserYanker.scala 47:17]
  wire [8:0] QueueCompatibility_31_io_deq_bits_tl_state_source; // @[UserYanker.scala 47:17]
  wire [4:0] QueueCompatibility_31_io_deq_bits_extra_id; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_31_io_covSum; // @[UserYanker.scala 47:17]
  wire  _ar_ready_WIRE_0 = QueueCompatibility_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _ar_ready_WIRE_1 = QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_1 = 4'h1 == auto_in_ar_bits_id ? _ar_ready_WIRE_1 : _ar_ready_WIRE_0; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_2 = QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_2 = 4'h2 == auto_in_ar_bits_id ? _ar_ready_WIRE_2 : _GEN_1; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_3 = QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_3 = 4'h3 == auto_in_ar_bits_id ? _ar_ready_WIRE_3 : _GEN_2; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_4 = QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_4 = 4'h4 == auto_in_ar_bits_id ? _ar_ready_WIRE_4 : _GEN_3; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_5 = QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_5 = 4'h5 == auto_in_ar_bits_id ? _ar_ready_WIRE_5 : _GEN_4; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_6 = QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_6 = 4'h6 == auto_in_ar_bits_id ? _ar_ready_WIRE_6 : _GEN_5; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_7 = QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_7 = 4'h7 == auto_in_ar_bits_id ? _ar_ready_WIRE_7 : _GEN_6; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_8 = QueueCompatibility_8_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_8 = 4'h8 == auto_in_ar_bits_id ? _ar_ready_WIRE_8 : _GEN_7; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_9 = QueueCompatibility_9_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_9 = 4'h9 == auto_in_ar_bits_id ? _ar_ready_WIRE_9 : _GEN_8; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_10 = QueueCompatibility_10_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_10 = 4'ha == auto_in_ar_bits_id ? _ar_ready_WIRE_10 : _GEN_9; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_11 = QueueCompatibility_11_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_11 = 4'hb == auto_in_ar_bits_id ? _ar_ready_WIRE_11 : _GEN_10; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_12 = QueueCompatibility_12_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_12 = 4'hc == auto_in_ar_bits_id ? _ar_ready_WIRE_12 : _GEN_11; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_13 = QueueCompatibility_13_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_13 = 4'hd == auto_in_ar_bits_id ? _ar_ready_WIRE_13 : _GEN_12; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_14 = QueueCompatibility_14_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_14 = 4'he == auto_in_ar_bits_id ? _ar_ready_WIRE_14 : _GEN_13; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_15 = QueueCompatibility_15_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_15 = 4'hf == auto_in_ar_bits_id ? _ar_ready_WIRE_15 : _GEN_14; // @[UserYanker.scala 56:{36,36}]
  wire  _r_valid_WIRE_0 = QueueCompatibility_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _r_valid_WIRE_1 = QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_17 = 4'h1 == auto_out_r_bits_id ? _r_valid_WIRE_1 : _r_valid_WIRE_0; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_2 = QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_18 = 4'h2 == auto_out_r_bits_id ? _r_valid_WIRE_2 : _GEN_17; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_3 = QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_19 = 4'h3 == auto_out_r_bits_id ? _r_valid_WIRE_3 : _GEN_18; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_4 = QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_20 = 4'h4 == auto_out_r_bits_id ? _r_valid_WIRE_4 : _GEN_19; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_5 = QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_21 = 4'h5 == auto_out_r_bits_id ? _r_valid_WIRE_5 : _GEN_20; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_6 = QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_22 = 4'h6 == auto_out_r_bits_id ? _r_valid_WIRE_6 : _GEN_21; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_7 = QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_23 = 4'h7 == auto_out_r_bits_id ? _r_valid_WIRE_7 : _GEN_22; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_8 = QueueCompatibility_8_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_24 = 4'h8 == auto_out_r_bits_id ? _r_valid_WIRE_8 : _GEN_23; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_9 = QueueCompatibility_9_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_25 = 4'h9 == auto_out_r_bits_id ? _r_valid_WIRE_9 : _GEN_24; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_10 = QueueCompatibility_10_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_26 = 4'ha == auto_out_r_bits_id ? _r_valid_WIRE_10 : _GEN_25; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_11 = QueueCompatibility_11_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_27 = 4'hb == auto_out_r_bits_id ? _r_valid_WIRE_11 : _GEN_26; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_12 = QueueCompatibility_12_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_28 = 4'hc == auto_out_r_bits_id ? _r_valid_WIRE_12 : _GEN_27; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_13 = QueueCompatibility_13_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_29 = 4'hd == auto_out_r_bits_id ? _r_valid_WIRE_13 : _GEN_28; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_14 = QueueCompatibility_14_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_30 = 4'he == auto_out_r_bits_id ? _r_valid_WIRE_14 : _GEN_29; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_15 = QueueCompatibility_15_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_31 = 4'hf == auto_out_r_bits_id ? _r_valid_WIRE_15 : _GEN_30; // @[UserYanker.scala 63:{28,28}]
  wire  _T_3 = ~reset; // @[UserYanker.scala 63:14]
  wire [4:0] _r_bits_WIRE_0_extra_id = QueueCompatibility_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _r_bits_WIRE_1_extra_id = QueueCompatibility_1_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_33 = 4'h1 == auto_out_r_bits_id ? _r_bits_WIRE_1_extra_id : _r_bits_WIRE_0_extra_id; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_2_extra_id = QueueCompatibility_2_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_34 = 4'h2 == auto_out_r_bits_id ? _r_bits_WIRE_2_extra_id : _GEN_33; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_3_extra_id = QueueCompatibility_3_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_35 = 4'h3 == auto_out_r_bits_id ? _r_bits_WIRE_3_extra_id : _GEN_34; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_4_extra_id = QueueCompatibility_4_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_36 = 4'h4 == auto_out_r_bits_id ? _r_bits_WIRE_4_extra_id : _GEN_35; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_5_extra_id = QueueCompatibility_5_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_37 = 4'h5 == auto_out_r_bits_id ? _r_bits_WIRE_5_extra_id : _GEN_36; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_6_extra_id = QueueCompatibility_6_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_38 = 4'h6 == auto_out_r_bits_id ? _r_bits_WIRE_6_extra_id : _GEN_37; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_7_extra_id = QueueCompatibility_7_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_39 = 4'h7 == auto_out_r_bits_id ? _r_bits_WIRE_7_extra_id : _GEN_38; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_8_extra_id = QueueCompatibility_8_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_40 = 4'h8 == auto_out_r_bits_id ? _r_bits_WIRE_8_extra_id : _GEN_39; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_9_extra_id = QueueCompatibility_9_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_41 = 4'h9 == auto_out_r_bits_id ? _r_bits_WIRE_9_extra_id : _GEN_40; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_10_extra_id = QueueCompatibility_10_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_42 = 4'ha == auto_out_r_bits_id ? _r_bits_WIRE_10_extra_id : _GEN_41; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_11_extra_id = QueueCompatibility_11_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_43 = 4'hb == auto_out_r_bits_id ? _r_bits_WIRE_11_extra_id : _GEN_42; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_12_extra_id = QueueCompatibility_12_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_44 = 4'hc == auto_out_r_bits_id ? _r_bits_WIRE_12_extra_id : _GEN_43; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_13_extra_id = QueueCompatibility_13_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_45 = 4'hd == auto_out_r_bits_id ? _r_bits_WIRE_13_extra_id : _GEN_44; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_14_extra_id = QueueCompatibility_14_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [4:0] _GEN_46 = 4'he == auto_out_r_bits_id ? _r_bits_WIRE_14_extra_id : _GEN_45; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _r_bits_WIRE_15_extra_id = QueueCompatibility_15_io_deq_bits_extra_id; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _r_bits_WIRE_0_tl_state_source = QueueCompatibility_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _r_bits_WIRE_1_tl_state_source = QueueCompatibility_1_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_49 = 4'h1 == auto_out_r_bits_id ? _r_bits_WIRE_1_tl_state_source : _r_bits_WIRE_0_tl_state_source; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_2_tl_state_source = QueueCompatibility_2_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_50 = 4'h2 == auto_out_r_bits_id ? _r_bits_WIRE_2_tl_state_source : _GEN_49; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_3_tl_state_source = QueueCompatibility_3_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_51 = 4'h3 == auto_out_r_bits_id ? _r_bits_WIRE_3_tl_state_source : _GEN_50; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_4_tl_state_source = QueueCompatibility_4_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_52 = 4'h4 == auto_out_r_bits_id ? _r_bits_WIRE_4_tl_state_source : _GEN_51; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_5_tl_state_source = QueueCompatibility_5_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_53 = 4'h5 == auto_out_r_bits_id ? _r_bits_WIRE_5_tl_state_source : _GEN_52; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_6_tl_state_source = QueueCompatibility_6_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_54 = 4'h6 == auto_out_r_bits_id ? _r_bits_WIRE_6_tl_state_source : _GEN_53; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_7_tl_state_source = QueueCompatibility_7_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_55 = 4'h7 == auto_out_r_bits_id ? _r_bits_WIRE_7_tl_state_source : _GEN_54; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_8_tl_state_source = QueueCompatibility_8_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_56 = 4'h8 == auto_out_r_bits_id ? _r_bits_WIRE_8_tl_state_source : _GEN_55; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_9_tl_state_source = QueueCompatibility_9_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_57 = 4'h9 == auto_out_r_bits_id ? _r_bits_WIRE_9_tl_state_source : _GEN_56; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_10_tl_state_source = QueueCompatibility_10_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_58 = 4'ha == auto_out_r_bits_id ? _r_bits_WIRE_10_tl_state_source : _GEN_57; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_11_tl_state_source = QueueCompatibility_11_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_59 = 4'hb == auto_out_r_bits_id ? _r_bits_WIRE_11_tl_state_source : _GEN_58; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_12_tl_state_source = QueueCompatibility_12_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_60 = 4'hc == auto_out_r_bits_id ? _r_bits_WIRE_12_tl_state_source : _GEN_59; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_13_tl_state_source = QueueCompatibility_13_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_61 = 4'hd == auto_out_r_bits_id ? _r_bits_WIRE_13_tl_state_source : _GEN_60; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_14_tl_state_source = QueueCompatibility_14_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [8:0] _GEN_62 = 4'he == auto_out_r_bits_id ? _r_bits_WIRE_14_tl_state_source : _GEN_61; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _r_bits_WIRE_15_tl_state_source = QueueCompatibility_15_io_deq_bits_tl_state_source; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _r_bits_WIRE_0_tl_state_size = QueueCompatibility_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _r_bits_WIRE_1_tl_state_size = QueueCompatibility_1_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_65 = 4'h1 == auto_out_r_bits_id ? _r_bits_WIRE_1_tl_state_size : _r_bits_WIRE_0_tl_state_size; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_2_tl_state_size = QueueCompatibility_2_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_66 = 4'h2 == auto_out_r_bits_id ? _r_bits_WIRE_2_tl_state_size : _GEN_65; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_3_tl_state_size = QueueCompatibility_3_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_67 = 4'h3 == auto_out_r_bits_id ? _r_bits_WIRE_3_tl_state_size : _GEN_66; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_4_tl_state_size = QueueCompatibility_4_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_68 = 4'h4 == auto_out_r_bits_id ? _r_bits_WIRE_4_tl_state_size : _GEN_67; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_5_tl_state_size = QueueCompatibility_5_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_69 = 4'h5 == auto_out_r_bits_id ? _r_bits_WIRE_5_tl_state_size : _GEN_68; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_6_tl_state_size = QueueCompatibility_6_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_70 = 4'h6 == auto_out_r_bits_id ? _r_bits_WIRE_6_tl_state_size : _GEN_69; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_7_tl_state_size = QueueCompatibility_7_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_71 = 4'h7 == auto_out_r_bits_id ? _r_bits_WIRE_7_tl_state_size : _GEN_70; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_8_tl_state_size = QueueCompatibility_8_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_72 = 4'h8 == auto_out_r_bits_id ? _r_bits_WIRE_8_tl_state_size : _GEN_71; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_9_tl_state_size = QueueCompatibility_9_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_73 = 4'h9 == auto_out_r_bits_id ? _r_bits_WIRE_9_tl_state_size : _GEN_72; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_10_tl_state_size = QueueCompatibility_10_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_74 = 4'ha == auto_out_r_bits_id ? _r_bits_WIRE_10_tl_state_size : _GEN_73; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_11_tl_state_size = QueueCompatibility_11_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_75 = 4'hb == auto_out_r_bits_id ? _r_bits_WIRE_11_tl_state_size : _GEN_74; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_12_tl_state_size = QueueCompatibility_12_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_76 = 4'hc == auto_out_r_bits_id ? _r_bits_WIRE_12_tl_state_size : _GEN_75; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_13_tl_state_size = QueueCompatibility_13_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_77 = 4'hd == auto_out_r_bits_id ? _r_bits_WIRE_13_tl_state_size : _GEN_76; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_14_tl_state_size = QueueCompatibility_14_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [3:0] _GEN_78 = 4'he == auto_out_r_bits_id ? _r_bits_WIRE_14_tl_state_size : _GEN_77; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _r_bits_WIRE_15_tl_state_size = QueueCompatibility_15_io_deq_bits_tl_state_size; // @[UserYanker.scala 62:{23,23}]
  wire [15:0] _arsel_T = 16'h1 << auto_in_ar_bits_id; // @[OneHot.scala 64:12]
  wire  arsel_0 = _arsel_T[0]; // @[UserYanker.scala 67:55]
  wire  arsel_1 = _arsel_T[1]; // @[UserYanker.scala 67:55]
  wire  arsel_2 = _arsel_T[2]; // @[UserYanker.scala 67:55]
  wire  arsel_3 = _arsel_T[3]; // @[UserYanker.scala 67:55]
  wire  arsel_4 = _arsel_T[4]; // @[UserYanker.scala 67:55]
  wire  arsel_5 = _arsel_T[5]; // @[UserYanker.scala 67:55]
  wire  arsel_6 = _arsel_T[6]; // @[UserYanker.scala 67:55]
  wire  arsel_7 = _arsel_T[7]; // @[UserYanker.scala 67:55]
  wire  arsel_8 = _arsel_T[8]; // @[UserYanker.scala 67:55]
  wire  arsel_9 = _arsel_T[9]; // @[UserYanker.scala 67:55]
  wire  arsel_10 = _arsel_T[10]; // @[UserYanker.scala 67:55]
  wire  arsel_11 = _arsel_T[11]; // @[UserYanker.scala 67:55]
  wire  arsel_12 = _arsel_T[12]; // @[UserYanker.scala 67:55]
  wire  arsel_13 = _arsel_T[13]; // @[UserYanker.scala 67:55]
  wire  arsel_14 = _arsel_T[14]; // @[UserYanker.scala 67:55]
  wire  arsel_15 = _arsel_T[15]; // @[UserYanker.scala 67:55]
  wire [15:0] _rsel_T = 16'h1 << auto_out_r_bits_id; // @[OneHot.scala 64:12]
  wire  rsel_0 = _rsel_T[0]; // @[UserYanker.scala 68:55]
  wire  rsel_1 = _rsel_T[1]; // @[UserYanker.scala 68:55]
  wire  rsel_2 = _rsel_T[2]; // @[UserYanker.scala 68:55]
  wire  rsel_3 = _rsel_T[3]; // @[UserYanker.scala 68:55]
  wire  rsel_4 = _rsel_T[4]; // @[UserYanker.scala 68:55]
  wire  rsel_5 = _rsel_T[5]; // @[UserYanker.scala 68:55]
  wire  rsel_6 = _rsel_T[6]; // @[UserYanker.scala 68:55]
  wire  rsel_7 = _rsel_T[7]; // @[UserYanker.scala 68:55]
  wire  rsel_8 = _rsel_T[8]; // @[UserYanker.scala 68:55]
  wire  rsel_9 = _rsel_T[9]; // @[UserYanker.scala 68:55]
  wire  rsel_10 = _rsel_T[10]; // @[UserYanker.scala 68:55]
  wire  rsel_11 = _rsel_T[11]; // @[UserYanker.scala 68:55]
  wire  rsel_12 = _rsel_T[12]; // @[UserYanker.scala 68:55]
  wire  rsel_13 = _rsel_T[13]; // @[UserYanker.scala 68:55]
  wire  rsel_14 = _rsel_T[14]; // @[UserYanker.scala 68:55]
  wire  rsel_15 = _rsel_T[15]; // @[UserYanker.scala 68:55]
  wire  _aw_ready_WIRE_0 = QueueCompatibility_16_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _aw_ready_WIRE_1 = QueueCompatibility_17_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_81 = 4'h1 == auto_in_aw_bits_id ? _aw_ready_WIRE_1 : _aw_ready_WIRE_0; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_2 = QueueCompatibility_18_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_82 = 4'h2 == auto_in_aw_bits_id ? _aw_ready_WIRE_2 : _GEN_81; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_3 = QueueCompatibility_19_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_83 = 4'h3 == auto_in_aw_bits_id ? _aw_ready_WIRE_3 : _GEN_82; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_4 = QueueCompatibility_20_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_84 = 4'h4 == auto_in_aw_bits_id ? _aw_ready_WIRE_4 : _GEN_83; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_5 = QueueCompatibility_21_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_85 = 4'h5 == auto_in_aw_bits_id ? _aw_ready_WIRE_5 : _GEN_84; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_6 = QueueCompatibility_22_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_86 = 4'h6 == auto_in_aw_bits_id ? _aw_ready_WIRE_6 : _GEN_85; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_7 = QueueCompatibility_23_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_87 = 4'h7 == auto_in_aw_bits_id ? _aw_ready_WIRE_7 : _GEN_86; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_8 = QueueCompatibility_24_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_88 = 4'h8 == auto_in_aw_bits_id ? _aw_ready_WIRE_8 : _GEN_87; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_9 = QueueCompatibility_25_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_89 = 4'h9 == auto_in_aw_bits_id ? _aw_ready_WIRE_9 : _GEN_88; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_10 = QueueCompatibility_26_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_90 = 4'ha == auto_in_aw_bits_id ? _aw_ready_WIRE_10 : _GEN_89; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_11 = QueueCompatibility_27_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_91 = 4'hb == auto_in_aw_bits_id ? _aw_ready_WIRE_11 : _GEN_90; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_12 = QueueCompatibility_28_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_92 = 4'hc == auto_in_aw_bits_id ? _aw_ready_WIRE_12 : _GEN_91; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_13 = QueueCompatibility_29_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_93 = 4'hd == auto_in_aw_bits_id ? _aw_ready_WIRE_13 : _GEN_92; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_14 = QueueCompatibility_30_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_94 = 4'he == auto_in_aw_bits_id ? _aw_ready_WIRE_14 : _GEN_93; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_15 = QueueCompatibility_31_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_95 = 4'hf == auto_in_aw_bits_id ? _aw_ready_WIRE_15 : _GEN_94; // @[UserYanker.scala 77:{36,36}]
  wire  _b_valid_WIRE_0 = QueueCompatibility_16_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _b_valid_WIRE_1 = QueueCompatibility_17_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_97 = 4'h1 == auto_out_b_bits_id ? _b_valid_WIRE_1 : _b_valid_WIRE_0; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_2 = QueueCompatibility_18_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_98 = 4'h2 == auto_out_b_bits_id ? _b_valid_WIRE_2 : _GEN_97; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_3 = QueueCompatibility_19_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_99 = 4'h3 == auto_out_b_bits_id ? _b_valid_WIRE_3 : _GEN_98; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_4 = QueueCompatibility_20_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_100 = 4'h4 == auto_out_b_bits_id ? _b_valid_WIRE_4 : _GEN_99; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_5 = QueueCompatibility_21_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_101 = 4'h5 == auto_out_b_bits_id ? _b_valid_WIRE_5 : _GEN_100; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_6 = QueueCompatibility_22_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_102 = 4'h6 == auto_out_b_bits_id ? _b_valid_WIRE_6 : _GEN_101; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_7 = QueueCompatibility_23_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_103 = 4'h7 == auto_out_b_bits_id ? _b_valid_WIRE_7 : _GEN_102; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_8 = QueueCompatibility_24_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_104 = 4'h8 == auto_out_b_bits_id ? _b_valid_WIRE_8 : _GEN_103; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_9 = QueueCompatibility_25_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_105 = 4'h9 == auto_out_b_bits_id ? _b_valid_WIRE_9 : _GEN_104; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_10 = QueueCompatibility_26_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_106 = 4'ha == auto_out_b_bits_id ? _b_valid_WIRE_10 : _GEN_105; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_11 = QueueCompatibility_27_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_107 = 4'hb == auto_out_b_bits_id ? _b_valid_WIRE_11 : _GEN_106; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_12 = QueueCompatibility_28_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_108 = 4'hc == auto_out_b_bits_id ? _b_valid_WIRE_12 : _GEN_107; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_13 = QueueCompatibility_29_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_109 = 4'hd == auto_out_b_bits_id ? _b_valid_WIRE_13 : _GEN_108; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_14 = QueueCompatibility_30_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_110 = 4'he == auto_out_b_bits_id ? _b_valid_WIRE_14 : _GEN_109; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_15 = QueueCompatibility_31_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_111 = 4'hf == auto_out_b_bits_id ? _b_valid_WIRE_15 : _GEN_110; // @[UserYanker.scala 84:{28,28}]
  wire [4:0] _b_bits_WIRE_0_extra_id = QueueCompatibility_16_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _b_bits_WIRE_1_extra_id = QueueCompatibility_17_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_113 = 4'h1 == auto_out_b_bits_id ? _b_bits_WIRE_1_extra_id : _b_bits_WIRE_0_extra_id; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_2_extra_id = QueueCompatibility_18_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_114 = 4'h2 == auto_out_b_bits_id ? _b_bits_WIRE_2_extra_id : _GEN_113; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_3_extra_id = QueueCompatibility_19_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_115 = 4'h3 == auto_out_b_bits_id ? _b_bits_WIRE_3_extra_id : _GEN_114; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_4_extra_id = QueueCompatibility_20_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_116 = 4'h4 == auto_out_b_bits_id ? _b_bits_WIRE_4_extra_id : _GEN_115; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_5_extra_id = QueueCompatibility_21_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_117 = 4'h5 == auto_out_b_bits_id ? _b_bits_WIRE_5_extra_id : _GEN_116; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_6_extra_id = QueueCompatibility_22_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_118 = 4'h6 == auto_out_b_bits_id ? _b_bits_WIRE_6_extra_id : _GEN_117; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_7_extra_id = QueueCompatibility_23_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_119 = 4'h7 == auto_out_b_bits_id ? _b_bits_WIRE_7_extra_id : _GEN_118; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_8_extra_id = QueueCompatibility_24_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_120 = 4'h8 == auto_out_b_bits_id ? _b_bits_WIRE_8_extra_id : _GEN_119; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_9_extra_id = QueueCompatibility_25_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_121 = 4'h9 == auto_out_b_bits_id ? _b_bits_WIRE_9_extra_id : _GEN_120; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_10_extra_id = QueueCompatibility_26_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_122 = 4'ha == auto_out_b_bits_id ? _b_bits_WIRE_10_extra_id : _GEN_121; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_11_extra_id = QueueCompatibility_27_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_123 = 4'hb == auto_out_b_bits_id ? _b_bits_WIRE_11_extra_id : _GEN_122; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_12_extra_id = QueueCompatibility_28_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_124 = 4'hc == auto_out_b_bits_id ? _b_bits_WIRE_12_extra_id : _GEN_123; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_13_extra_id = QueueCompatibility_29_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_125 = 4'hd == auto_out_b_bits_id ? _b_bits_WIRE_13_extra_id : _GEN_124; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_14_extra_id = QueueCompatibility_30_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [4:0] _GEN_126 = 4'he == auto_out_b_bits_id ? _b_bits_WIRE_14_extra_id : _GEN_125; // @[BundleMap.scala 247:{19,19}]
  wire [4:0] _b_bits_WIRE_15_extra_id = QueueCompatibility_31_io_deq_bits_extra_id; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _b_bits_WIRE_0_tl_state_source = QueueCompatibility_16_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _b_bits_WIRE_1_tl_state_source = QueueCompatibility_17_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_129 = 4'h1 == auto_out_b_bits_id ? _b_bits_WIRE_1_tl_state_source : _b_bits_WIRE_0_tl_state_source; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_2_tl_state_source = QueueCompatibility_18_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_130 = 4'h2 == auto_out_b_bits_id ? _b_bits_WIRE_2_tl_state_source : _GEN_129; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_3_tl_state_source = QueueCompatibility_19_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_131 = 4'h3 == auto_out_b_bits_id ? _b_bits_WIRE_3_tl_state_source : _GEN_130; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_4_tl_state_source = QueueCompatibility_20_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_132 = 4'h4 == auto_out_b_bits_id ? _b_bits_WIRE_4_tl_state_source : _GEN_131; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_5_tl_state_source = QueueCompatibility_21_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_133 = 4'h5 == auto_out_b_bits_id ? _b_bits_WIRE_5_tl_state_source : _GEN_132; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_6_tl_state_source = QueueCompatibility_22_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_134 = 4'h6 == auto_out_b_bits_id ? _b_bits_WIRE_6_tl_state_source : _GEN_133; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_7_tl_state_source = QueueCompatibility_23_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_135 = 4'h7 == auto_out_b_bits_id ? _b_bits_WIRE_7_tl_state_source : _GEN_134; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_8_tl_state_source = QueueCompatibility_24_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_136 = 4'h8 == auto_out_b_bits_id ? _b_bits_WIRE_8_tl_state_source : _GEN_135; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_9_tl_state_source = QueueCompatibility_25_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_137 = 4'h9 == auto_out_b_bits_id ? _b_bits_WIRE_9_tl_state_source : _GEN_136; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_10_tl_state_source = QueueCompatibility_26_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_138 = 4'ha == auto_out_b_bits_id ? _b_bits_WIRE_10_tl_state_source : _GEN_137; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_11_tl_state_source = QueueCompatibility_27_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_139 = 4'hb == auto_out_b_bits_id ? _b_bits_WIRE_11_tl_state_source : _GEN_138; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_12_tl_state_source = QueueCompatibility_28_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_140 = 4'hc == auto_out_b_bits_id ? _b_bits_WIRE_12_tl_state_source : _GEN_139; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_13_tl_state_source = QueueCompatibility_29_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_141 = 4'hd == auto_out_b_bits_id ? _b_bits_WIRE_13_tl_state_source : _GEN_140; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_14_tl_state_source = QueueCompatibility_30_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [8:0] _GEN_142 = 4'he == auto_out_b_bits_id ? _b_bits_WIRE_14_tl_state_source : _GEN_141; // @[BundleMap.scala 247:{19,19}]
  wire [8:0] _b_bits_WIRE_15_tl_state_source = QueueCompatibility_31_io_deq_bits_tl_state_source; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _b_bits_WIRE_0_tl_state_size = QueueCompatibility_16_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _b_bits_WIRE_1_tl_state_size = QueueCompatibility_17_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_145 = 4'h1 == auto_out_b_bits_id ? _b_bits_WIRE_1_tl_state_size : _b_bits_WIRE_0_tl_state_size; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_2_tl_state_size = QueueCompatibility_18_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_146 = 4'h2 == auto_out_b_bits_id ? _b_bits_WIRE_2_tl_state_size : _GEN_145; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_3_tl_state_size = QueueCompatibility_19_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_147 = 4'h3 == auto_out_b_bits_id ? _b_bits_WIRE_3_tl_state_size : _GEN_146; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_4_tl_state_size = QueueCompatibility_20_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_148 = 4'h4 == auto_out_b_bits_id ? _b_bits_WIRE_4_tl_state_size : _GEN_147; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_5_tl_state_size = QueueCompatibility_21_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_149 = 4'h5 == auto_out_b_bits_id ? _b_bits_WIRE_5_tl_state_size : _GEN_148; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_6_tl_state_size = QueueCompatibility_22_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_150 = 4'h6 == auto_out_b_bits_id ? _b_bits_WIRE_6_tl_state_size : _GEN_149; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_7_tl_state_size = QueueCompatibility_23_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_151 = 4'h7 == auto_out_b_bits_id ? _b_bits_WIRE_7_tl_state_size : _GEN_150; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_8_tl_state_size = QueueCompatibility_24_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_152 = 4'h8 == auto_out_b_bits_id ? _b_bits_WIRE_8_tl_state_size : _GEN_151; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_9_tl_state_size = QueueCompatibility_25_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_153 = 4'h9 == auto_out_b_bits_id ? _b_bits_WIRE_9_tl_state_size : _GEN_152; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_10_tl_state_size = QueueCompatibility_26_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_154 = 4'ha == auto_out_b_bits_id ? _b_bits_WIRE_10_tl_state_size : _GEN_153; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_11_tl_state_size = QueueCompatibility_27_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_155 = 4'hb == auto_out_b_bits_id ? _b_bits_WIRE_11_tl_state_size : _GEN_154; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_12_tl_state_size = QueueCompatibility_28_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_156 = 4'hc == auto_out_b_bits_id ? _b_bits_WIRE_12_tl_state_size : _GEN_155; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_13_tl_state_size = QueueCompatibility_29_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_157 = 4'hd == auto_out_b_bits_id ? _b_bits_WIRE_13_tl_state_size : _GEN_156; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_14_tl_state_size = QueueCompatibility_30_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [3:0] _GEN_158 = 4'he == auto_out_b_bits_id ? _b_bits_WIRE_14_tl_state_size : _GEN_157; // @[BundleMap.scala 247:{19,19}]
  wire [3:0] _b_bits_WIRE_15_tl_state_size = QueueCompatibility_31_io_deq_bits_tl_state_size; // @[UserYanker.scala 83:{23,23}]
  wire [15:0] _awsel_T = 16'h1 << auto_in_aw_bits_id; // @[OneHot.scala 64:12]
  wire  awsel_0 = _awsel_T[0]; // @[UserYanker.scala 88:55]
  wire  awsel_1 = _awsel_T[1]; // @[UserYanker.scala 88:55]
  wire  awsel_2 = _awsel_T[2]; // @[UserYanker.scala 88:55]
  wire  awsel_3 = _awsel_T[3]; // @[UserYanker.scala 88:55]
  wire  awsel_4 = _awsel_T[4]; // @[UserYanker.scala 88:55]
  wire  awsel_5 = _awsel_T[5]; // @[UserYanker.scala 88:55]
  wire  awsel_6 = _awsel_T[6]; // @[UserYanker.scala 88:55]
  wire  awsel_7 = _awsel_T[7]; // @[UserYanker.scala 88:55]
  wire  awsel_8 = _awsel_T[8]; // @[UserYanker.scala 88:55]
  wire  awsel_9 = _awsel_T[9]; // @[UserYanker.scala 88:55]
  wire  awsel_10 = _awsel_T[10]; // @[UserYanker.scala 88:55]
  wire  awsel_11 = _awsel_T[11]; // @[UserYanker.scala 88:55]
  wire  awsel_12 = _awsel_T[12]; // @[UserYanker.scala 88:55]
  wire  awsel_13 = _awsel_T[13]; // @[UserYanker.scala 88:55]
  wire  awsel_14 = _awsel_T[14]; // @[UserYanker.scala 88:55]
  wire  awsel_15 = _awsel_T[15]; // @[UserYanker.scala 88:55]
  wire [15:0] _bsel_T = 16'h1 << auto_out_b_bits_id; // @[OneHot.scala 64:12]
  wire  bsel_0 = _bsel_T[0]; // @[UserYanker.scala 89:55]
  wire  bsel_1 = _bsel_T[1]; // @[UserYanker.scala 89:55]
  wire  bsel_2 = _bsel_T[2]; // @[UserYanker.scala 89:55]
  wire  bsel_3 = _bsel_T[3]; // @[UserYanker.scala 89:55]
  wire  bsel_4 = _bsel_T[4]; // @[UserYanker.scala 89:55]
  wire  bsel_5 = _bsel_T[5]; // @[UserYanker.scala 89:55]
  wire  bsel_6 = _bsel_T[6]; // @[UserYanker.scala 89:55]
  wire  bsel_7 = _bsel_T[7]; // @[UserYanker.scala 89:55]
  wire  bsel_8 = _bsel_T[8]; // @[UserYanker.scala 89:55]
  wire  bsel_9 = _bsel_T[9]; // @[UserYanker.scala 89:55]
  wire  bsel_10 = _bsel_T[10]; // @[UserYanker.scala 89:55]
  wire  bsel_11 = _bsel_T[11]; // @[UserYanker.scala 89:55]
  wire  bsel_12 = _bsel_T[12]; // @[UserYanker.scala 89:55]
  wire  bsel_13 = _bsel_T[13]; // @[UserYanker.scala 89:55]
  wire  bsel_14 = _bsel_T[14]; // @[UserYanker.scala 89:55]
  wire  bsel_15 = _bsel_T[15]; // @[UserYanker.scala 89:55]
  wire [29:0] AXI4UserYanker_1_covSum;
  wire [29:0] QueueCompatibility_7_sum;
  wire [29:0] QueueCompatibility_30_sum;
  wire [29:0] QueueCompatibility_3_sum;
  wire [29:0] QueueCompatibility_31_sum;
  wire [29:0] QueueCompatibility_1_sum;
  wire [29:0] QueueCompatibility_19_sum;
  wire [29:0] QueueCompatibility_sum;
  wire [29:0] QueueCompatibility_27_sum;
  wire [29:0] QueueCompatibility_8_sum;
  wire [29:0] QueueCompatibility_29_sum;
  wire [29:0] QueueCompatibility_11_sum;
  wire [29:0] QueueCompatibility_21_sum;
  wire [29:0] QueueCompatibility_13_sum;
  wire [29:0] QueueCompatibility_14_sum;
  wire [29:0] QueueCompatibility_26_sum;
  wire [29:0] QueueCompatibility_24_sum;
  wire [29:0] QueueCompatibility_25_sum;
  wire [29:0] QueueCompatibility_16_sum;
  wire [29:0] QueueCompatibility_22_sum;
  wire [29:0] QueueCompatibility_12_sum;
  wire [29:0] QueueCompatibility_17_sum;
  wire [29:0] QueueCompatibility_28_sum;
  wire [29:0] QueueCompatibility_20_sum;
  wire [29:0] QueueCompatibility_18_sum;
  wire [29:0] QueueCompatibility_2_sum;
  wire [29:0] QueueCompatibility_4_sum;
  wire [29:0] QueueCompatibility_15_sum;
  wire [29:0] QueueCompatibility_6_sum;
  wire [29:0] QueueCompatibility_5_sum;
  wire [29:0] QueueCompatibility_23_sum;
  wire [29:0] QueueCompatibility_9_sum;
  wire [29:0] QueueCompatibility_10_sum;
  QueueCompatibility_4 QueueCompatibility ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_clock),
    .reset(QueueCompatibility_reset),
    .io_enq_ready(QueueCompatibility_io_enq_ready),
    .io_enq_valid(QueueCompatibility_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_io_deq_ready),
    .io_deq_valid(QueueCompatibility_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_1 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_1_clock),
    .reset(QueueCompatibility_1_reset),
    .io_enq_ready(QueueCompatibility_1_io_enq_ready),
    .io_enq_valid(QueueCompatibility_1_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_1_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_1_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_1_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_1_io_deq_ready),
    .io_deq_valid(QueueCompatibility_1_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_1_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_1_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_1_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_1_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_2 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_2_clock),
    .reset(QueueCompatibility_2_reset),
    .io_enq_ready(QueueCompatibility_2_io_enq_ready),
    .io_enq_valid(QueueCompatibility_2_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_2_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_2_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_2_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_2_io_deq_ready),
    .io_deq_valid(QueueCompatibility_2_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_2_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_2_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_2_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_2_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_3 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_3_clock),
    .reset(QueueCompatibility_3_reset),
    .io_enq_ready(QueueCompatibility_3_io_enq_ready),
    .io_enq_valid(QueueCompatibility_3_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_3_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_3_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_3_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_3_io_deq_ready),
    .io_deq_valid(QueueCompatibility_3_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_3_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_3_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_3_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_3_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_4 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_4_clock),
    .reset(QueueCompatibility_4_reset),
    .io_enq_ready(QueueCompatibility_4_io_enq_ready),
    .io_enq_valid(QueueCompatibility_4_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_4_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_4_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_4_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_4_io_deq_ready),
    .io_deq_valid(QueueCompatibility_4_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_4_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_4_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_4_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_4_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_5 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_5_clock),
    .reset(QueueCompatibility_5_reset),
    .io_enq_ready(QueueCompatibility_5_io_enq_ready),
    .io_enq_valid(QueueCompatibility_5_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_5_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_5_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_5_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_5_io_deq_ready),
    .io_deq_valid(QueueCompatibility_5_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_5_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_5_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_5_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_5_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_6 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_6_clock),
    .reset(QueueCompatibility_6_reset),
    .io_enq_ready(QueueCompatibility_6_io_enq_ready),
    .io_enq_valid(QueueCompatibility_6_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_6_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_6_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_6_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_6_io_deq_ready),
    .io_deq_valid(QueueCompatibility_6_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_6_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_6_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_6_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_6_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_7 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_7_clock),
    .reset(QueueCompatibility_7_reset),
    .io_enq_ready(QueueCompatibility_7_io_enq_ready),
    .io_enq_valid(QueueCompatibility_7_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_7_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_7_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_7_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_7_io_deq_ready),
    .io_deq_valid(QueueCompatibility_7_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_7_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_7_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_7_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_7_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_8 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_8_clock),
    .reset(QueueCompatibility_8_reset),
    .io_enq_ready(QueueCompatibility_8_io_enq_ready),
    .io_enq_valid(QueueCompatibility_8_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_8_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_8_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_8_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_8_io_deq_ready),
    .io_deq_valid(QueueCompatibility_8_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_8_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_8_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_8_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_8_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_9 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_9_clock),
    .reset(QueueCompatibility_9_reset),
    .io_enq_ready(QueueCompatibility_9_io_enq_ready),
    .io_enq_valid(QueueCompatibility_9_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_9_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_9_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_9_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_9_io_deq_ready),
    .io_deq_valid(QueueCompatibility_9_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_9_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_9_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_9_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_9_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_10 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_10_clock),
    .reset(QueueCompatibility_10_reset),
    .io_enq_ready(QueueCompatibility_10_io_enq_ready),
    .io_enq_valid(QueueCompatibility_10_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_10_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_10_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_10_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_10_io_deq_ready),
    .io_deq_valid(QueueCompatibility_10_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_10_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_10_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_10_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_10_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_11 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_11_clock),
    .reset(QueueCompatibility_11_reset),
    .io_enq_ready(QueueCompatibility_11_io_enq_ready),
    .io_enq_valid(QueueCompatibility_11_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_11_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_11_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_11_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_11_io_deq_ready),
    .io_deq_valid(QueueCompatibility_11_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_11_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_11_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_11_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_11_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_12 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_12_clock),
    .reset(QueueCompatibility_12_reset),
    .io_enq_ready(QueueCompatibility_12_io_enq_ready),
    .io_enq_valid(QueueCompatibility_12_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_12_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_12_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_12_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_12_io_deq_ready),
    .io_deq_valid(QueueCompatibility_12_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_12_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_12_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_12_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_12_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_13 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_13_clock),
    .reset(QueueCompatibility_13_reset),
    .io_enq_ready(QueueCompatibility_13_io_enq_ready),
    .io_enq_valid(QueueCompatibility_13_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_13_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_13_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_13_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_13_io_deq_ready),
    .io_deq_valid(QueueCompatibility_13_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_13_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_13_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_13_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_13_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_14 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_14_clock),
    .reset(QueueCompatibility_14_reset),
    .io_enq_ready(QueueCompatibility_14_io_enq_ready),
    .io_enq_valid(QueueCompatibility_14_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_14_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_14_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_14_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_14_io_deq_ready),
    .io_deq_valid(QueueCompatibility_14_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_14_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_14_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_14_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_14_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_15 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_15_clock),
    .reset(QueueCompatibility_15_reset),
    .io_enq_ready(QueueCompatibility_15_io_enq_ready),
    .io_enq_valid(QueueCompatibility_15_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_15_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_15_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_15_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_15_io_deq_ready),
    .io_deq_valid(QueueCompatibility_15_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_15_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_15_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_15_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_15_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_16 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_16_clock),
    .reset(QueueCompatibility_16_reset),
    .io_enq_ready(QueueCompatibility_16_io_enq_ready),
    .io_enq_valid(QueueCompatibility_16_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_16_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_16_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_16_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_16_io_deq_ready),
    .io_deq_valid(QueueCompatibility_16_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_16_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_16_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_16_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_16_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_17 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_17_clock),
    .reset(QueueCompatibility_17_reset),
    .io_enq_ready(QueueCompatibility_17_io_enq_ready),
    .io_enq_valid(QueueCompatibility_17_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_17_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_17_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_17_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_17_io_deq_ready),
    .io_deq_valid(QueueCompatibility_17_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_17_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_17_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_17_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_17_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_18 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_18_clock),
    .reset(QueueCompatibility_18_reset),
    .io_enq_ready(QueueCompatibility_18_io_enq_ready),
    .io_enq_valid(QueueCompatibility_18_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_18_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_18_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_18_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_18_io_deq_ready),
    .io_deq_valid(QueueCompatibility_18_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_18_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_18_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_18_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_18_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_19 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_19_clock),
    .reset(QueueCompatibility_19_reset),
    .io_enq_ready(QueueCompatibility_19_io_enq_ready),
    .io_enq_valid(QueueCompatibility_19_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_19_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_19_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_19_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_19_io_deq_ready),
    .io_deq_valid(QueueCompatibility_19_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_19_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_19_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_19_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_19_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_20 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_20_clock),
    .reset(QueueCompatibility_20_reset),
    .io_enq_ready(QueueCompatibility_20_io_enq_ready),
    .io_enq_valid(QueueCompatibility_20_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_20_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_20_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_20_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_20_io_deq_ready),
    .io_deq_valid(QueueCompatibility_20_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_20_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_20_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_20_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_20_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_21 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_21_clock),
    .reset(QueueCompatibility_21_reset),
    .io_enq_ready(QueueCompatibility_21_io_enq_ready),
    .io_enq_valid(QueueCompatibility_21_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_21_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_21_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_21_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_21_io_deq_ready),
    .io_deq_valid(QueueCompatibility_21_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_21_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_21_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_21_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_21_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_22 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_22_clock),
    .reset(QueueCompatibility_22_reset),
    .io_enq_ready(QueueCompatibility_22_io_enq_ready),
    .io_enq_valid(QueueCompatibility_22_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_22_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_22_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_22_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_22_io_deq_ready),
    .io_deq_valid(QueueCompatibility_22_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_22_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_22_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_22_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_22_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_23 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_23_clock),
    .reset(QueueCompatibility_23_reset),
    .io_enq_ready(QueueCompatibility_23_io_enq_ready),
    .io_enq_valid(QueueCompatibility_23_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_23_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_23_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_23_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_23_io_deq_ready),
    .io_deq_valid(QueueCompatibility_23_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_23_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_23_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_23_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_23_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_24 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_24_clock),
    .reset(QueueCompatibility_24_reset),
    .io_enq_ready(QueueCompatibility_24_io_enq_ready),
    .io_enq_valid(QueueCompatibility_24_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_24_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_24_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_24_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_24_io_deq_ready),
    .io_deq_valid(QueueCompatibility_24_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_24_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_24_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_24_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_24_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_25 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_25_clock),
    .reset(QueueCompatibility_25_reset),
    .io_enq_ready(QueueCompatibility_25_io_enq_ready),
    .io_enq_valid(QueueCompatibility_25_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_25_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_25_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_25_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_25_io_deq_ready),
    .io_deq_valid(QueueCompatibility_25_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_25_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_25_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_25_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_25_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_26 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_26_clock),
    .reset(QueueCompatibility_26_reset),
    .io_enq_ready(QueueCompatibility_26_io_enq_ready),
    .io_enq_valid(QueueCompatibility_26_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_26_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_26_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_26_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_26_io_deq_ready),
    .io_deq_valid(QueueCompatibility_26_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_26_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_26_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_26_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_26_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_27 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_27_clock),
    .reset(QueueCompatibility_27_reset),
    .io_enq_ready(QueueCompatibility_27_io_enq_ready),
    .io_enq_valid(QueueCompatibility_27_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_27_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_27_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_27_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_27_io_deq_ready),
    .io_deq_valid(QueueCompatibility_27_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_27_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_27_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_27_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_27_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_28 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_28_clock),
    .reset(QueueCompatibility_28_reset),
    .io_enq_ready(QueueCompatibility_28_io_enq_ready),
    .io_enq_valid(QueueCompatibility_28_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_28_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_28_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_28_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_28_io_deq_ready),
    .io_deq_valid(QueueCompatibility_28_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_28_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_28_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_28_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_28_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_29 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_29_clock),
    .reset(QueueCompatibility_29_reset),
    .io_enq_ready(QueueCompatibility_29_io_enq_ready),
    .io_enq_valid(QueueCompatibility_29_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_29_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_29_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_29_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_29_io_deq_ready),
    .io_deq_valid(QueueCompatibility_29_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_29_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_29_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_29_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_29_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_30 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_30_clock),
    .reset(QueueCompatibility_30_reset),
    .io_enq_ready(QueueCompatibility_30_io_enq_ready),
    .io_enq_valid(QueueCompatibility_30_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_30_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_30_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_30_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_30_io_deq_ready),
    .io_deq_valid(QueueCompatibility_30_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_30_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_30_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_30_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_30_io_covSum)
  );
  QueueCompatibility_4 QueueCompatibility_31 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_31_clock),
    .reset(QueueCompatibility_31_reset),
    .io_enq_ready(QueueCompatibility_31_io_enq_ready),
    .io_enq_valid(QueueCompatibility_31_io_enq_valid),
    .io_enq_bits_tl_state_size(QueueCompatibility_31_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(QueueCompatibility_31_io_enq_bits_tl_state_source),
    .io_enq_bits_extra_id(QueueCompatibility_31_io_enq_bits_extra_id),
    .io_deq_ready(QueueCompatibility_31_io_deq_ready),
    .io_deq_valid(QueueCompatibility_31_io_deq_valid),
    .io_deq_bits_tl_state_size(QueueCompatibility_31_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(QueueCompatibility_31_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id(QueueCompatibility_31_io_deq_bits_extra_id),
    .io_covSum(QueueCompatibility_31_io_covSum)
  );
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_95; // @[UserYanker.scala 77:36]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_echo_tl_state_size = 4'hf == auto_out_b_bits_id ? _b_bits_WIRE_15_tl_state_size : _GEN_158; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_b_bits_echo_tl_state_source = 4'hf == auto_out_b_bits_id ? _b_bits_WIRE_15_tl_state_source : _GEN_142; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_b_bits_echo_extra_id = 4'hf == auto_out_b_bits_id ? _b_bits_WIRE_15_extra_id : _GEN_126; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_15; // @[UserYanker.scala 56:36]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_echo_tl_state_size = 4'hf == auto_out_r_bits_id ? _r_bits_WIRE_15_tl_state_size : _GEN_78; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_echo_tl_state_source = 4'hf == auto_out_r_bits_id ? _r_bits_WIRE_15_tl_state_source : _GEN_62; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_echo_extra_id = 4'hf == auto_out_r_bits_id ? _r_bits_WIRE_15_extra_id : _GEN_46; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_95; // @[UserYanker.scala 78:36]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_valid = auto_in_w_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_15; // @[UserYanker.scala 57:36]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_clock = clock;
  assign QueueCompatibility_reset = reset;
  assign QueueCompatibility_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_0; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_0 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_1_clock = clock;
  assign QueueCompatibility_1_reset = reset;
  assign QueueCompatibility_1_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_1; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_1_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_1 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_2_clock = clock;
  assign QueueCompatibility_2_reset = reset;
  assign QueueCompatibility_2_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_2; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_2_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_2 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_3_clock = clock;
  assign QueueCompatibility_3_reset = reset;
  assign QueueCompatibility_3_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_3; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_3_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_3 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_4_clock = clock;
  assign QueueCompatibility_4_reset = reset;
  assign QueueCompatibility_4_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_4; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_4_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_4_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_4_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_4_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_4 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_5_clock = clock;
  assign QueueCompatibility_5_reset = reset;
  assign QueueCompatibility_5_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_5; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_5_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_5_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_5_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_5_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_5 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_6_clock = clock;
  assign QueueCompatibility_6_reset = reset;
  assign QueueCompatibility_6_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_6; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_6_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_6_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_6_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_6_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_6 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_7_clock = clock;
  assign QueueCompatibility_7_reset = reset;
  assign QueueCompatibility_7_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_7; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_7_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_7_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_7_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_7_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_7 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_8_clock = clock;
  assign QueueCompatibility_8_reset = reset;
  assign QueueCompatibility_8_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_8; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_8_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_8_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_8_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_8_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_8 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_9_clock = clock;
  assign QueueCompatibility_9_reset = reset;
  assign QueueCompatibility_9_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_9; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_9_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_9_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_9_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_9_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_9 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_10_clock = clock;
  assign QueueCompatibility_10_reset = reset;
  assign QueueCompatibility_10_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_10; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_10_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_10_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_10_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_10_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_10 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_11_clock = clock;
  assign QueueCompatibility_11_reset = reset;
  assign QueueCompatibility_11_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_11; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_11_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_11_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_11_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_11_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_11 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_12_clock = clock;
  assign QueueCompatibility_12_reset = reset;
  assign QueueCompatibility_12_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_12; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_12_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_12_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_12_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_12_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_12 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_13_clock = clock;
  assign QueueCompatibility_13_reset = reset;
  assign QueueCompatibility_13_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_13; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_13_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_13_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_13_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_13_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_13 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_14_clock = clock;
  assign QueueCompatibility_14_reset = reset;
  assign QueueCompatibility_14_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_14; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_14_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_14_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_14_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_14_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_14 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_15_clock = clock;
  assign QueueCompatibility_15_reset = reset;
  assign QueueCompatibility_15_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_15; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_15_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_15_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_15_io_enq_bits_extra_id = auto_in_ar_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_15_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_15 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_16_clock = clock;
  assign QueueCompatibility_16_reset = reset;
  assign QueueCompatibility_16_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_0; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_16_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_16_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_16_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_16_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_0; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_17_clock = clock;
  assign QueueCompatibility_17_reset = reset;
  assign QueueCompatibility_17_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_1; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_17_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_17_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_17_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_17_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_1; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_18_clock = clock;
  assign QueueCompatibility_18_reset = reset;
  assign QueueCompatibility_18_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_2; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_18_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_18_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_18_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_18_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_2; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_19_clock = clock;
  assign QueueCompatibility_19_reset = reset;
  assign QueueCompatibility_19_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_3; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_19_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_19_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_19_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_19_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_3; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_20_clock = clock;
  assign QueueCompatibility_20_reset = reset;
  assign QueueCompatibility_20_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_4; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_20_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_20_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_20_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_20_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_4; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_21_clock = clock;
  assign QueueCompatibility_21_reset = reset;
  assign QueueCompatibility_21_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_5; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_21_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_21_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_21_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_21_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_5; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_22_clock = clock;
  assign QueueCompatibility_22_reset = reset;
  assign QueueCompatibility_22_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_6; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_22_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_22_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_22_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_22_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_6; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_23_clock = clock;
  assign QueueCompatibility_23_reset = reset;
  assign QueueCompatibility_23_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_7; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_23_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_23_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_23_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_23_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_7; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_24_clock = clock;
  assign QueueCompatibility_24_reset = reset;
  assign QueueCompatibility_24_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_8; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_24_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_24_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_24_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_24_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_8; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_25_clock = clock;
  assign QueueCompatibility_25_reset = reset;
  assign QueueCompatibility_25_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_9; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_25_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_25_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_25_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_25_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_9; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_26_clock = clock;
  assign QueueCompatibility_26_reset = reset;
  assign QueueCompatibility_26_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_10; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_26_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_26_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_26_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_26_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_10; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_27_clock = clock;
  assign QueueCompatibility_27_reset = reset;
  assign QueueCompatibility_27_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_11; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_27_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_27_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_27_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_27_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_11; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_28_clock = clock;
  assign QueueCompatibility_28_reset = reset;
  assign QueueCompatibility_28_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_12; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_28_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_28_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_28_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_28_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_12; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_29_clock = clock;
  assign QueueCompatibility_29_reset = reset;
  assign QueueCompatibility_29_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_13; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_29_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_29_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_29_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_29_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_13; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_30_clock = clock;
  assign QueueCompatibility_30_reset = reset;
  assign QueueCompatibility_30_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_14; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_30_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_30_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_30_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_30_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_14; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_31_clock = clock;
  assign QueueCompatibility_31_reset = reset;
  assign QueueCompatibility_31_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_15; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_31_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_31_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_31_io_enq_bits_extra_id = auto_in_aw_bits_echo_extra_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_31_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_15; // @[UserYanker.scala 91:53]
  assign AXI4UserYanker_1_covSum = 30'h0;
  assign QueueCompatibility_7_sum = AXI4UserYanker_1_covSum + QueueCompatibility_7_io_covSum;
  assign QueueCompatibility_30_sum = QueueCompatibility_7_sum + QueueCompatibility_30_io_covSum;
  assign QueueCompatibility_3_sum = QueueCompatibility_30_sum + QueueCompatibility_3_io_covSum;
  assign QueueCompatibility_31_sum = QueueCompatibility_3_sum + QueueCompatibility_31_io_covSum;
  assign QueueCompatibility_1_sum = QueueCompatibility_31_sum + QueueCompatibility_1_io_covSum;
  assign QueueCompatibility_19_sum = QueueCompatibility_1_sum + QueueCompatibility_19_io_covSum;
  assign QueueCompatibility_sum = QueueCompatibility_19_sum + QueueCompatibility_io_covSum;
  assign QueueCompatibility_27_sum = QueueCompatibility_sum + QueueCompatibility_27_io_covSum;
  assign QueueCompatibility_8_sum = QueueCompatibility_27_sum + QueueCompatibility_8_io_covSum;
  assign QueueCompatibility_29_sum = QueueCompatibility_8_sum + QueueCompatibility_29_io_covSum;
  assign QueueCompatibility_11_sum = QueueCompatibility_29_sum + QueueCompatibility_11_io_covSum;
  assign QueueCompatibility_21_sum = QueueCompatibility_11_sum + QueueCompatibility_21_io_covSum;
  assign QueueCompatibility_13_sum = QueueCompatibility_21_sum + QueueCompatibility_13_io_covSum;
  assign QueueCompatibility_14_sum = QueueCompatibility_13_sum + QueueCompatibility_14_io_covSum;
  assign QueueCompatibility_26_sum = QueueCompatibility_14_sum + QueueCompatibility_26_io_covSum;
  assign QueueCompatibility_24_sum = QueueCompatibility_26_sum + QueueCompatibility_24_io_covSum;
  assign QueueCompatibility_25_sum = QueueCompatibility_24_sum + QueueCompatibility_25_io_covSum;
  assign QueueCompatibility_16_sum = QueueCompatibility_25_sum + QueueCompatibility_16_io_covSum;
  assign QueueCompatibility_22_sum = QueueCompatibility_16_sum + QueueCompatibility_22_io_covSum;
  assign QueueCompatibility_12_sum = QueueCompatibility_22_sum + QueueCompatibility_12_io_covSum;
  assign QueueCompatibility_17_sum = QueueCompatibility_12_sum + QueueCompatibility_17_io_covSum;
  assign QueueCompatibility_28_sum = QueueCompatibility_17_sum + QueueCompatibility_28_io_covSum;
  assign QueueCompatibility_20_sum = QueueCompatibility_28_sum + QueueCompatibility_20_io_covSum;
  assign QueueCompatibility_18_sum = QueueCompatibility_20_sum + QueueCompatibility_18_io_covSum;
  assign QueueCompatibility_2_sum = QueueCompatibility_18_sum + QueueCompatibility_2_io_covSum;
  assign QueueCompatibility_4_sum = QueueCompatibility_2_sum + QueueCompatibility_4_io_covSum;
  assign QueueCompatibility_15_sum = QueueCompatibility_4_sum + QueueCompatibility_15_io_covSum;
  assign QueueCompatibility_6_sum = QueueCompatibility_15_sum + QueueCompatibility_6_io_covSum;
  assign QueueCompatibility_5_sum = QueueCompatibility_6_sum + QueueCompatibility_5_io_covSum;
  assign QueueCompatibility_23_sum = QueueCompatibility_5_sum + QueueCompatibility_23_io_covSum;
  assign QueueCompatibility_9_sum = QueueCompatibility_23_sum + QueueCompatibility_9_io_covSum;
  assign QueueCompatibility_10_sum = QueueCompatibility_9_sum + QueueCompatibility_10_io_covSum;
  assign io_covSum = QueueCompatibility_10_sum;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_r_valid | _GEN_31) & ~reset) begin
          $fatal; // @[UserYanker.scala 63:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_out_r_valid | _GEN_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:63 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 63:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_b_valid | _GEN_111) & _T_3) begin
          $fatal; // @[UserYanker.scala 84:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~auto_out_b_valid | _GEN_111)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:84 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 84:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4IdIndexer_1(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [8:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
  input  [3:0]  auto_in_aw_bits_echo_tl_state_size,
  input  [8:0]  auto_in_aw_bits_echo_tl_state_source,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [8:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [3:0]  auto_in_b_bits_echo_tl_state_size,
  output [8:0]  auto_in_b_bits_echo_tl_state_source,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [8:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
  input  [3:0]  auto_in_ar_bits_echo_tl_state_size,
  input  [8:0]  auto_in_ar_bits_echo_tl_state_source,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [8:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [3:0]  auto_in_r_bits_echo_tl_state_size,
  output [8:0]  auto_in_r_bits_echo_tl_state_source,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  output [3:0]  auto_out_aw_bits_echo_tl_state_size,
  output [8:0]  auto_out_aw_bits_echo_tl_state_source,
  output [4:0]  auto_out_aw_bits_echo_extra_id,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [3:0]  auto_out_b_bits_echo_tl_state_size,
  input  [8:0]  auto_out_b_bits_echo_tl_state_source,
  input  [4:0]  auto_out_b_bits_echo_extra_id,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output [3:0]  auto_out_ar_bits_echo_tl_state_size,
  output [8:0]  auto_out_ar_bits_echo_tl_state_source,
  output [4:0]  auto_out_ar_bits_echo_extra_id,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [3:0]  auto_out_r_bits_echo_tl_state_size,
  input  [8:0]  auto_out_r_bits_echo_tl_state_source,
  input  [4:0]  auto_out_r_bits_echo_extra_id,
  input         auto_out_r_bits_last,
  output [29:0] io_covSum
);
  wire [29:0] AXI4IdIndexer_1_covSum;
  assign auto_in_aw_ready = auto_out_aw_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_id = {auto_out_b_bits_echo_extra_id,auto_out_b_bits_id}; // @[Cat.scala 31:58]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_echo_tl_state_size = auto_out_b_bits_echo_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_echo_tl_state_source = auto_out_b_bits_echo_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_id = {auto_out_r_bits_echo_extra_id,auto_out_r_bits_id}; // @[Cat.scala 31:58]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_echo_tl_state_size = auto_out_r_bits_echo_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id[3:0]; // @[Nodes.scala 1207:84 BundleMap.scala 247:19]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_echo_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_echo_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_echo_extra_id = auto_in_aw_bits_id[8:4]; // @[IdIndexer.scala 71:56]
  assign auto_out_w_valid = auto_in_w_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id[3:0]; // @[Nodes.scala 1207:84 BundleMap.scala 247:19]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_echo_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_echo_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_echo_extra_id = auto_in_ar_bits_id[8:4]; // @[IdIndexer.scala 70:56]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign AXI4IdIndexer_1_covSum = 30'h0;
  assign io_covSum = AXI4IdIndexer_1_covSum;
endmodule
module Queue_19(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [8:0]  io_enq_bits_id,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_cache,
  input  [2:0]  io_enq_bits_prot,
  input  [3:0]  io_enq_bits_echo_tl_state_size,
  input  [8:0]  io_enq_bits_echo_tl_state_source,
  input         io_enq_bits_wen,
  input         io_deq_ready,
  output        io_deq_valid,
  output [8:0]  io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output        io_deq_bits_lock,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [3:0]  io_deq_bits_qos,
  output [3:0]  io_deq_bits_echo_tl_state_size,
  output [8:0]  io_deq_bits_echo_tl_state_source,
  output        io_deq_bits_wen,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] ram_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [8:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [8:0] ram_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_len [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_burst [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_lock [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_lock_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_lock_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_lock_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_lock_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_lock_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_lock_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_cache [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_cache_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_cache_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_cache_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_prot [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_prot_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_prot_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_prot_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_qos [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_qos_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_qos_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_qos_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_qos_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_qos_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_qos_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_echo_tl_state_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_echo_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_echo_tl_state_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [8:0] ram_echo_tl_state_source [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [8:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [8:0] ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_wen [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_wen_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_wen_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wen_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wen_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_wen_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_wen_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_wen_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_20 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_20 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  reg  Queue_19_covState; // @[Register tracking Queue_19 state]
  reg  Queue_19_covMap [0:1]; // @[Coverage map for Queue_19]
  wire  Queue_19_covMap_read_en; // @[Coverage map for Queue_19]
  wire  Queue_19_covMap_read_addr; // @[Coverage map for Queue_19]
  wire  Queue_19_covMap_read_data; // @[Coverage map for Queue_19]
  wire  Queue_19_covMap_write_data; // @[Coverage map for Queue_19]
  wire  Queue_19_covMap_write_addr; // @[Coverage map for Queue_19]
  wire  Queue_19_covMap_write_mask; // @[Coverage map for Queue_19]
  wire  Queue_19_covMap_write_en; // @[Coverage map for Queue_19]
  reg [29:0] Queue_19_covSum; // @[Sum of coverage map]
  wire  maybe_full_shl;
  wire  maybe_full_pad;
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_burst_MPORT_data = 2'h1;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_lock_io_deq_bits_MPORT_en = 1'h1;
  assign ram_lock_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_lock_io_deq_bits_MPORT_data = ram_lock[ram_lock_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_lock_MPORT_data = 1'h0;
  assign ram_lock_MPORT_addr = 1'h0;
  assign ram_lock_MPORT_mask = 1'h1;
  assign ram_lock_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_cache_io_deq_bits_MPORT_en = 1'h1;
  assign ram_cache_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_cache_io_deq_bits_MPORT_data = ram_cache[ram_cache_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_cache_MPORT_data = io_enq_bits_cache;
  assign ram_cache_MPORT_addr = 1'h0;
  assign ram_cache_MPORT_mask = 1'h1;
  assign ram_cache_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_prot_io_deq_bits_MPORT_en = 1'h1;
  assign ram_prot_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_prot_io_deq_bits_MPORT_data = ram_prot[ram_prot_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_prot_MPORT_data = io_enq_bits_prot;
  assign ram_prot_MPORT_addr = 1'h0;
  assign ram_prot_MPORT_mask = 1'h1;
  assign ram_prot_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_qos_io_deq_bits_MPORT_en = 1'h1;
  assign ram_qos_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_qos_io_deq_bits_MPORT_data = ram_qos[ram_qos_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_qos_MPORT_data = 4'h0;
  assign ram_qos_MPORT_addr = 1'h0;
  assign ram_qos_MPORT_mask = 1'h1;
  assign ram_qos_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_echo_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_size_io_deq_bits_MPORT_data =
    ram_echo_tl_state_size[ram_echo_tl_state_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_echo_tl_state_size_MPORT_data = io_enq_bits_echo_tl_state_size;
  assign ram_echo_tl_state_size_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_size_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_size_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign ram_wen_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wen_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wen_io_deq_bits_MPORT_data = ram_wen[ram_wen_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_wen_MPORT_data = io_enq_bits_wen;
  assign ram_wen_MPORT_addr = 1'h0;
  assign ram_wen_MPORT_mask = 1'h1;
  assign ram_wen_MPORT_en = empty ? _GEN_20 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_burst = empty ? 2'h1 : ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_lock = empty ? 1'h0 : ram_lock_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_cache = empty ? io_enq_bits_cache : ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_prot = empty ? io_enq_bits_prot : ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_qos = empty ? 4'h0 : ram_qos_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_echo_tl_state_size = empty ? io_enq_bits_echo_tl_state_size :
    ram_echo_tl_state_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_echo_tl_state_source = empty ? io_enq_bits_echo_tl_state_source :
    ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_wen = empty ? io_enq_bits_wen : ram_wen_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign Queue_19_covMap_read_en = 1'h1;
  assign Queue_19_covMap_read_addr = Queue_19_covState;
  assign Queue_19_covMap_read_data = Queue_19_covMap[Queue_19_covMap_read_addr]; // @[Coverage map for Queue_19]
  assign Queue_19_covMap_write_data = 1'h1;
  assign Queue_19_covMap_write_addr = Queue_19_covState;
  assign Queue_19_covMap_write_mask = 1'h1;
  assign Queue_19_covMap_write_en = ~metaReset;
  assign maybe_full_shl = maybe_full;
  assign maybe_full_pad = maybe_full_shl;
  assign io_covSum = Queue_19_covSum;
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_lock_MPORT_en & ram_lock_MPORT_mask) begin
      ram_lock[ram_lock_MPORT_addr] <= ram_lock_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_cache_MPORT_en & ram_cache_MPORT_mask) begin
      ram_cache[ram_cache_MPORT_addr] <= ram_cache_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_prot_MPORT_en & ram_prot_MPORT_mask) begin
      ram_prot[ram_prot_MPORT_addr] <= ram_prot_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_qos_MPORT_en & ram_qos_MPORT_mask) begin
      ram_qos[ram_qos_MPORT_addr] <= ram_qos_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_echo_tl_state_size_MPORT_en & ram_echo_tl_state_size_MPORT_mask) begin
      ram_echo_tl_state_size[ram_echo_tl_state_size_MPORT_addr] <= ram_echo_tl_state_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_wen_MPORT_en & ram_wen_MPORT_mask) begin
      ram_wen[ram_wen_MPORT_addr] <= ram_wen_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
    Queue_19_covState <= maybe_full_pad;
    if (Queue_19_covMap_write_en & Queue_19_covMap_write_mask) begin
      Queue_19_covMap[Queue_19_covMap_write_addr] <= Queue_19_covMap_write_data; // @[Coverage map for Queue_19]
    end
    if (!(Queue_19_covMap_read_data | metaReset)) begin
      Queue_19_covSum <= Queue_19_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_lock[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_qos[initvar] = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_echo_tl_state_size[initvar] = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_echo_tl_state_source[initvar] = _RAND_10[8:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wen[initvar] = _RAND_11[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Queue_19_covMap[initvar] = 0; //_14[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  maybe_full = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  Queue_19_covState = 0; //_13[0:0];
  _RAND_15 = {1{`RANDOM}};
  Queue_19_covSum = 0; //_15[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLToAXI4(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [8:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input         auto_in_a_bits_user_amba_prot_bufferable,
  input         auto_in_a_bits_user_amba_prot_modifiable,
  input         auto_in_a_bits_user_amba_prot_readalloc,
  input         auto_in_a_bits_user_amba_prot_writealloc,
  input         auto_in_a_bits_user_amba_prot_privileged,
  input         auto_in_a_bits_user_amba_prot_secure,
  input         auto_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [8:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [8:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  output [3:0]  auto_out_aw_bits_echo_tl_state_size,
  output [8:0]  auto_out_aw_bits_echo_tl_state_source,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [8:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input  [3:0]  auto_out_b_bits_echo_tl_state_size,
  input  [8:0]  auto_out_b_bits_echo_tl_state_source,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [8:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output [3:0]  auto_out_ar_bits_echo_tl_state_size,
  output [8:0]  auto_out_ar_bits_echo_tl_state_source,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [8:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input  [3:0]  auto_out_r_bits_echo_tl_state_size,
  input  [8:0]  auto_out_r_bits_echo_tl_state_source,
  input         auto_out_r_bits_last,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_519;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_520;
`endif // RANDOMIZE_REG_INIT
  wire  deq_clock; // @[Decoupled.scala 361:21]
  wire  deq_reset; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [63:0] deq_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] deq_io_enq_bits_strb; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_bits_last; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [63:0] deq_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] deq_io_deq_bits_strb; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_bits_last; // @[Decoupled.scala 361:21]
  wire [29:0] deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  deq_metaReset; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_clock; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_reset; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [8:0] queue_arw_deq_io_enq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] queue_arw_deq_io_enq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] queue_arw_deq_io_enq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] queue_arw_deq_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] queue_arw_deq_io_enq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] queue_arw_deq_io_enq_bits_prot; // @[Decoupled.scala 361:21]
  wire [3:0] queue_arw_deq_io_enq_bits_echo_tl_state_size; // @[Decoupled.scala 361:21]
  wire [8:0] queue_arw_deq_io_enq_bits_echo_tl_state_source; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_io_enq_bits_wen; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [8:0] queue_arw_deq_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] queue_arw_deq_io_deq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] queue_arw_deq_io_deq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] queue_arw_deq_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] queue_arw_deq_io_deq_bits_burst; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_io_deq_bits_lock; // @[Decoupled.scala 361:21]
  wire [3:0] queue_arw_deq_io_deq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] queue_arw_deq_io_deq_bits_prot; // @[Decoupled.scala 361:21]
  wire [3:0] queue_arw_deq_io_deq_bits_qos; // @[Decoupled.scala 361:21]
  wire [3:0] queue_arw_deq_io_deq_bits_echo_tl_state_size; // @[Decoupled.scala 361:21]
  wire [8:0] queue_arw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_io_deq_bits_wen; // @[Decoupled.scala 361:21]
  wire [29:0] queue_arw_deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  queue_arw_deq_metaReset; // @[Decoupled.scala 361:21]
  wire  a_isPut = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  reg  count_512; // @[ToAXI4.scala 254:28]
  wire  idle_511 = ~count_512; // @[ToAXI4.scala 256:26]
  reg  count_511; // @[ToAXI4.scala 254:28]
  wire  idle_510 = ~count_511; // @[ToAXI4.scala 256:26]
  reg  count_510; // @[ToAXI4.scala 254:28]
  wire  idle_509 = ~count_510; // @[ToAXI4.scala 256:26]
  reg  count_509; // @[ToAXI4.scala 254:28]
  wire  idle_508 = ~count_509; // @[ToAXI4.scala 256:26]
  reg  count_508; // @[ToAXI4.scala 254:28]
  wire  idle_507 = ~count_508; // @[ToAXI4.scala 256:26]
  reg  count_507; // @[ToAXI4.scala 254:28]
  wire  idle_506 = ~count_507; // @[ToAXI4.scala 256:26]
  reg  count_506; // @[ToAXI4.scala 254:28]
  wire  idle_505 = ~count_506; // @[ToAXI4.scala 256:26]
  reg  count_505; // @[ToAXI4.scala 254:28]
  wire  idle_504 = ~count_505; // @[ToAXI4.scala 256:26]
  reg  count_504; // @[ToAXI4.scala 254:28]
  wire  idle_503 = ~count_504; // @[ToAXI4.scala 256:26]
  reg  count_503; // @[ToAXI4.scala 254:28]
  wire  idle_502 = ~count_503; // @[ToAXI4.scala 256:26]
  reg  count_502; // @[ToAXI4.scala 254:28]
  wire  idle_501 = ~count_502; // @[ToAXI4.scala 256:26]
  reg  count_501; // @[ToAXI4.scala 254:28]
  wire  idle_500 = ~count_501; // @[ToAXI4.scala 256:26]
  reg  count_500; // @[ToAXI4.scala 254:28]
  wire  idle_499 = ~count_500; // @[ToAXI4.scala 256:26]
  reg  count_499; // @[ToAXI4.scala 254:28]
  wire  idle_498 = ~count_499; // @[ToAXI4.scala 256:26]
  reg  count_498; // @[ToAXI4.scala 254:28]
  wire  idle_497 = ~count_498; // @[ToAXI4.scala 256:26]
  reg  count_497; // @[ToAXI4.scala 254:28]
  wire  idle_496 = ~count_497; // @[ToAXI4.scala 256:26]
  reg  count_496; // @[ToAXI4.scala 254:28]
  wire  idle_495 = ~count_496; // @[ToAXI4.scala 256:26]
  reg  count_495; // @[ToAXI4.scala 254:28]
  wire  idle_494 = ~count_495; // @[ToAXI4.scala 256:26]
  reg  count_494; // @[ToAXI4.scala 254:28]
  wire  idle_493 = ~count_494; // @[ToAXI4.scala 256:26]
  reg  count_493; // @[ToAXI4.scala 254:28]
  wire  idle_492 = ~count_493; // @[ToAXI4.scala 256:26]
  reg  count_492; // @[ToAXI4.scala 254:28]
  wire  idle_491 = ~count_492; // @[ToAXI4.scala 256:26]
  reg  count_491; // @[ToAXI4.scala 254:28]
  wire  idle_490 = ~count_491; // @[ToAXI4.scala 256:26]
  reg  count_490; // @[ToAXI4.scala 254:28]
  wire  idle_489 = ~count_490; // @[ToAXI4.scala 256:26]
  reg  count_489; // @[ToAXI4.scala 254:28]
  wire  idle_488 = ~count_489; // @[ToAXI4.scala 256:26]
  reg  count_488; // @[ToAXI4.scala 254:28]
  wire  idle_487 = ~count_488; // @[ToAXI4.scala 256:26]
  reg  count_487; // @[ToAXI4.scala 254:28]
  wire  idle_486 = ~count_487; // @[ToAXI4.scala 256:26]
  reg  count_486; // @[ToAXI4.scala 254:28]
  wire  idle_485 = ~count_486; // @[ToAXI4.scala 256:26]
  reg  count_485; // @[ToAXI4.scala 254:28]
  wire  idle_484 = ~count_485; // @[ToAXI4.scala 256:26]
  reg  count_484; // @[ToAXI4.scala 254:28]
  wire  idle_483 = ~count_484; // @[ToAXI4.scala 256:26]
  reg  count_483; // @[ToAXI4.scala 254:28]
  wire  idle_482 = ~count_483; // @[ToAXI4.scala 256:26]
  reg  count_482; // @[ToAXI4.scala 254:28]
  wire  idle_481 = ~count_482; // @[ToAXI4.scala 256:26]
  reg  count_481; // @[ToAXI4.scala 254:28]
  wire  idle_480 = ~count_481; // @[ToAXI4.scala 256:26]
  reg  count_480; // @[ToAXI4.scala 254:28]
  wire  idle_479 = ~count_480; // @[ToAXI4.scala 256:26]
  reg  count_479; // @[ToAXI4.scala 254:28]
  wire  idle_478 = ~count_479; // @[ToAXI4.scala 256:26]
  reg  count_478; // @[ToAXI4.scala 254:28]
  wire  idle_477 = ~count_478; // @[ToAXI4.scala 256:26]
  reg  count_477; // @[ToAXI4.scala 254:28]
  wire  idle_476 = ~count_477; // @[ToAXI4.scala 256:26]
  reg  count_476; // @[ToAXI4.scala 254:28]
  wire  idle_475 = ~count_476; // @[ToAXI4.scala 256:26]
  reg  count_475; // @[ToAXI4.scala 254:28]
  wire  idle_474 = ~count_475; // @[ToAXI4.scala 256:26]
  reg  count_474; // @[ToAXI4.scala 254:28]
  wire  idle_473 = ~count_474; // @[ToAXI4.scala 256:26]
  reg  count_473; // @[ToAXI4.scala 254:28]
  wire  idle_472 = ~count_473; // @[ToAXI4.scala 256:26]
  reg  count_472; // @[ToAXI4.scala 254:28]
  wire  idle_471 = ~count_472; // @[ToAXI4.scala 256:26]
  reg  count_471; // @[ToAXI4.scala 254:28]
  wire  idle_470 = ~count_471; // @[ToAXI4.scala 256:26]
  reg  count_470; // @[ToAXI4.scala 254:28]
  wire  idle_469 = ~count_470; // @[ToAXI4.scala 256:26]
  reg  count_469; // @[ToAXI4.scala 254:28]
  wire  idle_468 = ~count_469; // @[ToAXI4.scala 256:26]
  reg  count_468; // @[ToAXI4.scala 254:28]
  wire  idle_467 = ~count_468; // @[ToAXI4.scala 256:26]
  reg  count_467; // @[ToAXI4.scala 254:28]
  wire  idle_466 = ~count_467; // @[ToAXI4.scala 256:26]
  reg  count_466; // @[ToAXI4.scala 254:28]
  wire  idle_465 = ~count_466; // @[ToAXI4.scala 256:26]
  reg  count_465; // @[ToAXI4.scala 254:28]
  wire  idle_464 = ~count_465; // @[ToAXI4.scala 256:26]
  reg  count_464; // @[ToAXI4.scala 254:28]
  wire  idle_463 = ~count_464; // @[ToAXI4.scala 256:26]
  reg  count_463; // @[ToAXI4.scala 254:28]
  wire  idle_462 = ~count_463; // @[ToAXI4.scala 256:26]
  reg  count_462; // @[ToAXI4.scala 254:28]
  wire  idle_461 = ~count_462; // @[ToAXI4.scala 256:26]
  reg  count_461; // @[ToAXI4.scala 254:28]
  wire  idle_460 = ~count_461; // @[ToAXI4.scala 256:26]
  reg  count_460; // @[ToAXI4.scala 254:28]
  wire  idle_459 = ~count_460; // @[ToAXI4.scala 256:26]
  reg  count_459; // @[ToAXI4.scala 254:28]
  wire  idle_458 = ~count_459; // @[ToAXI4.scala 256:26]
  reg  count_458; // @[ToAXI4.scala 254:28]
  wire  idle_457 = ~count_458; // @[ToAXI4.scala 256:26]
  reg  count_457; // @[ToAXI4.scala 254:28]
  wire  idle_456 = ~count_457; // @[ToAXI4.scala 256:26]
  reg  count_456; // @[ToAXI4.scala 254:28]
  wire  idle_455 = ~count_456; // @[ToAXI4.scala 256:26]
  reg  count_455; // @[ToAXI4.scala 254:28]
  wire  idle_454 = ~count_455; // @[ToAXI4.scala 256:26]
  reg  count_454; // @[ToAXI4.scala 254:28]
  wire  idle_453 = ~count_454; // @[ToAXI4.scala 256:26]
  reg  count_453; // @[ToAXI4.scala 254:28]
  wire  idle_452 = ~count_453; // @[ToAXI4.scala 256:26]
  reg  count_452; // @[ToAXI4.scala 254:28]
  wire  idle_451 = ~count_452; // @[ToAXI4.scala 256:26]
  reg  count_451; // @[ToAXI4.scala 254:28]
  wire  idle_450 = ~count_451; // @[ToAXI4.scala 256:26]
  reg  count_450; // @[ToAXI4.scala 254:28]
  wire  idle_449 = ~count_450; // @[ToAXI4.scala 256:26]
  reg  count_449; // @[ToAXI4.scala 254:28]
  wire  idle_448 = ~count_449; // @[ToAXI4.scala 256:26]
  reg  count_448; // @[ToAXI4.scala 254:28]
  wire  idle_447 = ~count_448; // @[ToAXI4.scala 256:26]
  reg  count_447; // @[ToAXI4.scala 254:28]
  wire  idle_446 = ~count_447; // @[ToAXI4.scala 256:26]
  reg  count_446; // @[ToAXI4.scala 254:28]
  wire  idle_445 = ~count_446; // @[ToAXI4.scala 256:26]
  reg  count_445; // @[ToAXI4.scala 254:28]
  wire  idle_444 = ~count_445; // @[ToAXI4.scala 256:26]
  reg  count_444; // @[ToAXI4.scala 254:28]
  wire  idle_443 = ~count_444; // @[ToAXI4.scala 256:26]
  reg  count_443; // @[ToAXI4.scala 254:28]
  wire  idle_442 = ~count_443; // @[ToAXI4.scala 256:26]
  reg  count_442; // @[ToAXI4.scala 254:28]
  wire  idle_441 = ~count_442; // @[ToAXI4.scala 256:26]
  reg  count_441; // @[ToAXI4.scala 254:28]
  wire  idle_440 = ~count_441; // @[ToAXI4.scala 256:26]
  reg  count_440; // @[ToAXI4.scala 254:28]
  wire  idle_439 = ~count_440; // @[ToAXI4.scala 256:26]
  reg  count_439; // @[ToAXI4.scala 254:28]
  wire  idle_438 = ~count_439; // @[ToAXI4.scala 256:26]
  reg  count_438; // @[ToAXI4.scala 254:28]
  wire  idle_437 = ~count_438; // @[ToAXI4.scala 256:26]
  reg  count_437; // @[ToAXI4.scala 254:28]
  wire  idle_436 = ~count_437; // @[ToAXI4.scala 256:26]
  reg  count_436; // @[ToAXI4.scala 254:28]
  wire  idle_435 = ~count_436; // @[ToAXI4.scala 256:26]
  reg  count_435; // @[ToAXI4.scala 254:28]
  wire  idle_434 = ~count_435; // @[ToAXI4.scala 256:26]
  reg  count_434; // @[ToAXI4.scala 254:28]
  wire  idle_433 = ~count_434; // @[ToAXI4.scala 256:26]
  reg  count_433; // @[ToAXI4.scala 254:28]
  wire  idle_432 = ~count_433; // @[ToAXI4.scala 256:26]
  reg  count_432; // @[ToAXI4.scala 254:28]
  wire  idle_431 = ~count_432; // @[ToAXI4.scala 256:26]
  reg  count_431; // @[ToAXI4.scala 254:28]
  wire  idle_430 = ~count_431; // @[ToAXI4.scala 256:26]
  reg  count_430; // @[ToAXI4.scala 254:28]
  wire  idle_429 = ~count_430; // @[ToAXI4.scala 256:26]
  reg  count_429; // @[ToAXI4.scala 254:28]
  wire  idle_428 = ~count_429; // @[ToAXI4.scala 256:26]
  reg  count_428; // @[ToAXI4.scala 254:28]
  wire  idle_427 = ~count_428; // @[ToAXI4.scala 256:26]
  reg  count_427; // @[ToAXI4.scala 254:28]
  wire  idle_426 = ~count_427; // @[ToAXI4.scala 256:26]
  reg  count_426; // @[ToAXI4.scala 254:28]
  wire  idle_425 = ~count_426; // @[ToAXI4.scala 256:26]
  reg  count_425; // @[ToAXI4.scala 254:28]
  wire  idle_424 = ~count_425; // @[ToAXI4.scala 256:26]
  reg  count_424; // @[ToAXI4.scala 254:28]
  wire  idle_423 = ~count_424; // @[ToAXI4.scala 256:26]
  reg  count_423; // @[ToAXI4.scala 254:28]
  wire  idle_422 = ~count_423; // @[ToAXI4.scala 256:26]
  reg  count_422; // @[ToAXI4.scala 254:28]
  wire  idle_421 = ~count_422; // @[ToAXI4.scala 256:26]
  reg  count_421; // @[ToAXI4.scala 254:28]
  wire  idle_420 = ~count_421; // @[ToAXI4.scala 256:26]
  reg  count_420; // @[ToAXI4.scala 254:28]
  wire  idle_419 = ~count_420; // @[ToAXI4.scala 256:26]
  reg  count_419; // @[ToAXI4.scala 254:28]
  wire  idle_418 = ~count_419; // @[ToAXI4.scala 256:26]
  reg  count_418; // @[ToAXI4.scala 254:28]
  wire  idle_417 = ~count_418; // @[ToAXI4.scala 256:26]
  reg  count_417; // @[ToAXI4.scala 254:28]
  wire  idle_416 = ~count_417; // @[ToAXI4.scala 256:26]
  reg  count_416; // @[ToAXI4.scala 254:28]
  wire  idle_415 = ~count_416; // @[ToAXI4.scala 256:26]
  reg  count_415; // @[ToAXI4.scala 254:28]
  wire  idle_414 = ~count_415; // @[ToAXI4.scala 256:26]
  reg  count_414; // @[ToAXI4.scala 254:28]
  wire  idle_413 = ~count_414; // @[ToAXI4.scala 256:26]
  reg  count_413; // @[ToAXI4.scala 254:28]
  wire  idle_412 = ~count_413; // @[ToAXI4.scala 256:26]
  reg  count_412; // @[ToAXI4.scala 254:28]
  wire  idle_411 = ~count_412; // @[ToAXI4.scala 256:26]
  reg  count_411; // @[ToAXI4.scala 254:28]
  wire  idle_410 = ~count_411; // @[ToAXI4.scala 256:26]
  reg  count_410; // @[ToAXI4.scala 254:28]
  wire  idle_409 = ~count_410; // @[ToAXI4.scala 256:26]
  reg  count_409; // @[ToAXI4.scala 254:28]
  wire  idle_408 = ~count_409; // @[ToAXI4.scala 256:26]
  reg  count_408; // @[ToAXI4.scala 254:28]
  wire  idle_407 = ~count_408; // @[ToAXI4.scala 256:26]
  reg  count_407; // @[ToAXI4.scala 254:28]
  wire  idle_406 = ~count_407; // @[ToAXI4.scala 256:26]
  reg  count_406; // @[ToAXI4.scala 254:28]
  wire  idle_405 = ~count_406; // @[ToAXI4.scala 256:26]
  reg  count_405; // @[ToAXI4.scala 254:28]
  wire  idle_404 = ~count_405; // @[ToAXI4.scala 256:26]
  reg  count_404; // @[ToAXI4.scala 254:28]
  wire  idle_403 = ~count_404; // @[ToAXI4.scala 256:26]
  reg  count_403; // @[ToAXI4.scala 254:28]
  wire  idle_402 = ~count_403; // @[ToAXI4.scala 256:26]
  reg  count_402; // @[ToAXI4.scala 254:28]
  wire  idle_401 = ~count_402; // @[ToAXI4.scala 256:26]
  reg  count_401; // @[ToAXI4.scala 254:28]
  wire  idle_400 = ~count_401; // @[ToAXI4.scala 256:26]
  reg  count_400; // @[ToAXI4.scala 254:28]
  wire  idle_399 = ~count_400; // @[ToAXI4.scala 256:26]
  reg  count_399; // @[ToAXI4.scala 254:28]
  wire  idle_398 = ~count_399; // @[ToAXI4.scala 256:26]
  reg  count_398; // @[ToAXI4.scala 254:28]
  wire  idle_397 = ~count_398; // @[ToAXI4.scala 256:26]
  reg  count_397; // @[ToAXI4.scala 254:28]
  wire  idle_396 = ~count_397; // @[ToAXI4.scala 256:26]
  reg  count_396; // @[ToAXI4.scala 254:28]
  wire  idle_395 = ~count_396; // @[ToAXI4.scala 256:26]
  reg  count_395; // @[ToAXI4.scala 254:28]
  wire  idle_394 = ~count_395; // @[ToAXI4.scala 256:26]
  reg  count_394; // @[ToAXI4.scala 254:28]
  wire  idle_393 = ~count_394; // @[ToAXI4.scala 256:26]
  reg  count_393; // @[ToAXI4.scala 254:28]
  wire  idle_392 = ~count_393; // @[ToAXI4.scala 256:26]
  reg  count_392; // @[ToAXI4.scala 254:28]
  wire  idle_391 = ~count_392; // @[ToAXI4.scala 256:26]
  reg  count_391; // @[ToAXI4.scala 254:28]
  wire  idle_390 = ~count_391; // @[ToAXI4.scala 256:26]
  reg  count_390; // @[ToAXI4.scala 254:28]
  wire  idle_389 = ~count_390; // @[ToAXI4.scala 256:26]
  reg  count_389; // @[ToAXI4.scala 254:28]
  wire  idle_388 = ~count_389; // @[ToAXI4.scala 256:26]
  reg  count_388; // @[ToAXI4.scala 254:28]
  wire  idle_387 = ~count_388; // @[ToAXI4.scala 256:26]
  reg  count_387; // @[ToAXI4.scala 254:28]
  wire  idle_386 = ~count_387; // @[ToAXI4.scala 256:26]
  reg  count_386; // @[ToAXI4.scala 254:28]
  wire  idle_385 = ~count_386; // @[ToAXI4.scala 256:26]
  reg  count_385; // @[ToAXI4.scala 254:28]
  wire  idle_384 = ~count_385; // @[ToAXI4.scala 256:26]
  reg  count_384; // @[ToAXI4.scala 254:28]
  wire  idle_383 = ~count_384; // @[ToAXI4.scala 256:26]
  reg  count_383; // @[ToAXI4.scala 254:28]
  wire  idle_382 = ~count_383; // @[ToAXI4.scala 256:26]
  reg  count_382; // @[ToAXI4.scala 254:28]
  wire  idle_381 = ~count_382; // @[ToAXI4.scala 256:26]
  reg  count_381; // @[ToAXI4.scala 254:28]
  wire  idle_380 = ~count_381; // @[ToAXI4.scala 256:26]
  reg  count_380; // @[ToAXI4.scala 254:28]
  wire  idle_379 = ~count_380; // @[ToAXI4.scala 256:26]
  reg  count_379; // @[ToAXI4.scala 254:28]
  wire  idle_378 = ~count_379; // @[ToAXI4.scala 256:26]
  reg  count_378; // @[ToAXI4.scala 254:28]
  wire  idle_377 = ~count_378; // @[ToAXI4.scala 256:26]
  reg  count_377; // @[ToAXI4.scala 254:28]
  wire  idle_376 = ~count_377; // @[ToAXI4.scala 256:26]
  reg  count_376; // @[ToAXI4.scala 254:28]
  wire  idle_375 = ~count_376; // @[ToAXI4.scala 256:26]
  reg  count_375; // @[ToAXI4.scala 254:28]
  wire  idle_374 = ~count_375; // @[ToAXI4.scala 256:26]
  reg  count_374; // @[ToAXI4.scala 254:28]
  wire  idle_373 = ~count_374; // @[ToAXI4.scala 256:26]
  reg  count_373; // @[ToAXI4.scala 254:28]
  wire  idle_372 = ~count_373; // @[ToAXI4.scala 256:26]
  reg  count_372; // @[ToAXI4.scala 254:28]
  wire  idle_371 = ~count_372; // @[ToAXI4.scala 256:26]
  reg  count_371; // @[ToAXI4.scala 254:28]
  wire  idle_370 = ~count_371; // @[ToAXI4.scala 256:26]
  reg  count_370; // @[ToAXI4.scala 254:28]
  wire  idle_369 = ~count_370; // @[ToAXI4.scala 256:26]
  reg  count_369; // @[ToAXI4.scala 254:28]
  wire  idle_368 = ~count_369; // @[ToAXI4.scala 256:26]
  reg  count_368; // @[ToAXI4.scala 254:28]
  wire  idle_367 = ~count_368; // @[ToAXI4.scala 256:26]
  reg  count_367; // @[ToAXI4.scala 254:28]
  wire  idle_366 = ~count_367; // @[ToAXI4.scala 256:26]
  reg  count_366; // @[ToAXI4.scala 254:28]
  wire  idle_365 = ~count_366; // @[ToAXI4.scala 256:26]
  reg  count_365; // @[ToAXI4.scala 254:28]
  wire  idle_364 = ~count_365; // @[ToAXI4.scala 256:26]
  reg  count_364; // @[ToAXI4.scala 254:28]
  wire  idle_363 = ~count_364; // @[ToAXI4.scala 256:26]
  reg  count_363; // @[ToAXI4.scala 254:28]
  wire  idle_362 = ~count_363; // @[ToAXI4.scala 256:26]
  reg  count_362; // @[ToAXI4.scala 254:28]
  wire  idle_361 = ~count_362; // @[ToAXI4.scala 256:26]
  reg  count_361; // @[ToAXI4.scala 254:28]
  wire  idle_360 = ~count_361; // @[ToAXI4.scala 256:26]
  reg  count_360; // @[ToAXI4.scala 254:28]
  wire  idle_359 = ~count_360; // @[ToAXI4.scala 256:26]
  reg  count_359; // @[ToAXI4.scala 254:28]
  wire  idle_358 = ~count_359; // @[ToAXI4.scala 256:26]
  reg  count_358; // @[ToAXI4.scala 254:28]
  wire  idle_357 = ~count_358; // @[ToAXI4.scala 256:26]
  reg  count_357; // @[ToAXI4.scala 254:28]
  wire  idle_356 = ~count_357; // @[ToAXI4.scala 256:26]
  reg  count_356; // @[ToAXI4.scala 254:28]
  wire  idle_355 = ~count_356; // @[ToAXI4.scala 256:26]
  reg  count_355; // @[ToAXI4.scala 254:28]
  wire  idle_354 = ~count_355; // @[ToAXI4.scala 256:26]
  reg  count_354; // @[ToAXI4.scala 254:28]
  wire  idle_353 = ~count_354; // @[ToAXI4.scala 256:26]
  reg  count_353; // @[ToAXI4.scala 254:28]
  wire  idle_352 = ~count_353; // @[ToAXI4.scala 256:26]
  reg  count_352; // @[ToAXI4.scala 254:28]
  wire  idle_351 = ~count_352; // @[ToAXI4.scala 256:26]
  reg  count_351; // @[ToAXI4.scala 254:28]
  wire  idle_350 = ~count_351; // @[ToAXI4.scala 256:26]
  reg  count_350; // @[ToAXI4.scala 254:28]
  wire  idle_349 = ~count_350; // @[ToAXI4.scala 256:26]
  reg  count_349; // @[ToAXI4.scala 254:28]
  wire  idle_348 = ~count_349; // @[ToAXI4.scala 256:26]
  reg  count_348; // @[ToAXI4.scala 254:28]
  wire  idle_347 = ~count_348; // @[ToAXI4.scala 256:26]
  reg  count_347; // @[ToAXI4.scala 254:28]
  wire  idle_346 = ~count_347; // @[ToAXI4.scala 256:26]
  reg  count_346; // @[ToAXI4.scala 254:28]
  wire  idle_345 = ~count_346; // @[ToAXI4.scala 256:26]
  reg  count_345; // @[ToAXI4.scala 254:28]
  wire  idle_344 = ~count_345; // @[ToAXI4.scala 256:26]
  reg  count_344; // @[ToAXI4.scala 254:28]
  wire  idle_343 = ~count_344; // @[ToAXI4.scala 256:26]
  reg  count_343; // @[ToAXI4.scala 254:28]
  wire  idle_342 = ~count_343; // @[ToAXI4.scala 256:26]
  reg  count_342; // @[ToAXI4.scala 254:28]
  wire  idle_341 = ~count_342; // @[ToAXI4.scala 256:26]
  reg  count_341; // @[ToAXI4.scala 254:28]
  wire  idle_340 = ~count_341; // @[ToAXI4.scala 256:26]
  reg  count_340; // @[ToAXI4.scala 254:28]
  wire  idle_339 = ~count_340; // @[ToAXI4.scala 256:26]
  reg  count_339; // @[ToAXI4.scala 254:28]
  wire  idle_338 = ~count_339; // @[ToAXI4.scala 256:26]
  reg  count_338; // @[ToAXI4.scala 254:28]
  wire  idle_337 = ~count_338; // @[ToAXI4.scala 256:26]
  reg  count_337; // @[ToAXI4.scala 254:28]
  wire  idle_336 = ~count_337; // @[ToAXI4.scala 256:26]
  reg  count_336; // @[ToAXI4.scala 254:28]
  wire  idle_335 = ~count_336; // @[ToAXI4.scala 256:26]
  reg  count_335; // @[ToAXI4.scala 254:28]
  wire  idle_334 = ~count_335; // @[ToAXI4.scala 256:26]
  reg  count_334; // @[ToAXI4.scala 254:28]
  wire  idle_333 = ~count_334; // @[ToAXI4.scala 256:26]
  reg  count_333; // @[ToAXI4.scala 254:28]
  wire  idle_332 = ~count_333; // @[ToAXI4.scala 256:26]
  reg  count_332; // @[ToAXI4.scala 254:28]
  wire  idle_331 = ~count_332; // @[ToAXI4.scala 256:26]
  reg  count_331; // @[ToAXI4.scala 254:28]
  wire  idle_330 = ~count_331; // @[ToAXI4.scala 256:26]
  reg  count_330; // @[ToAXI4.scala 254:28]
  wire  idle_329 = ~count_330; // @[ToAXI4.scala 256:26]
  reg  count_329; // @[ToAXI4.scala 254:28]
  wire  idle_328 = ~count_329; // @[ToAXI4.scala 256:26]
  reg  count_328; // @[ToAXI4.scala 254:28]
  wire  idle_327 = ~count_328; // @[ToAXI4.scala 256:26]
  reg  count_327; // @[ToAXI4.scala 254:28]
  wire  idle_326 = ~count_327; // @[ToAXI4.scala 256:26]
  reg  count_326; // @[ToAXI4.scala 254:28]
  wire  idle_325 = ~count_326; // @[ToAXI4.scala 256:26]
  reg  count_325; // @[ToAXI4.scala 254:28]
  wire  idle_324 = ~count_325; // @[ToAXI4.scala 256:26]
  reg  count_324; // @[ToAXI4.scala 254:28]
  wire  idle_323 = ~count_324; // @[ToAXI4.scala 256:26]
  reg  count_323; // @[ToAXI4.scala 254:28]
  wire  idle_322 = ~count_323; // @[ToAXI4.scala 256:26]
  reg  count_322; // @[ToAXI4.scala 254:28]
  wire  idle_321 = ~count_322; // @[ToAXI4.scala 256:26]
  reg  count_321; // @[ToAXI4.scala 254:28]
  wire  idle_320 = ~count_321; // @[ToAXI4.scala 256:26]
  reg  count_320; // @[ToAXI4.scala 254:28]
  wire  idle_319 = ~count_320; // @[ToAXI4.scala 256:26]
  reg  count_319; // @[ToAXI4.scala 254:28]
  wire  idle_318 = ~count_319; // @[ToAXI4.scala 256:26]
  reg  count_318; // @[ToAXI4.scala 254:28]
  wire  idle_317 = ~count_318; // @[ToAXI4.scala 256:26]
  reg  count_317; // @[ToAXI4.scala 254:28]
  wire  idle_316 = ~count_317; // @[ToAXI4.scala 256:26]
  reg  count_316; // @[ToAXI4.scala 254:28]
  wire  idle_315 = ~count_316; // @[ToAXI4.scala 256:26]
  reg  count_315; // @[ToAXI4.scala 254:28]
  wire  idle_314 = ~count_315; // @[ToAXI4.scala 256:26]
  reg  count_314; // @[ToAXI4.scala 254:28]
  wire  idle_313 = ~count_314; // @[ToAXI4.scala 256:26]
  reg  count_313; // @[ToAXI4.scala 254:28]
  wire  idle_312 = ~count_313; // @[ToAXI4.scala 256:26]
  reg  count_312; // @[ToAXI4.scala 254:28]
  wire  idle_311 = ~count_312; // @[ToAXI4.scala 256:26]
  reg  count_311; // @[ToAXI4.scala 254:28]
  wire  idle_310 = ~count_311; // @[ToAXI4.scala 256:26]
  reg  count_310; // @[ToAXI4.scala 254:28]
  wire  idle_309 = ~count_310; // @[ToAXI4.scala 256:26]
  reg  count_309; // @[ToAXI4.scala 254:28]
  wire  idle_308 = ~count_309; // @[ToAXI4.scala 256:26]
  reg  count_308; // @[ToAXI4.scala 254:28]
  wire  idle_307 = ~count_308; // @[ToAXI4.scala 256:26]
  reg  count_307; // @[ToAXI4.scala 254:28]
  wire  idle_306 = ~count_307; // @[ToAXI4.scala 256:26]
  reg  count_306; // @[ToAXI4.scala 254:28]
  wire  idle_305 = ~count_306; // @[ToAXI4.scala 256:26]
  reg  count_305; // @[ToAXI4.scala 254:28]
  wire  idle_304 = ~count_305; // @[ToAXI4.scala 256:26]
  reg  count_304; // @[ToAXI4.scala 254:28]
  wire  idle_303 = ~count_304; // @[ToAXI4.scala 256:26]
  reg  count_303; // @[ToAXI4.scala 254:28]
  wire  idle_302 = ~count_303; // @[ToAXI4.scala 256:26]
  reg  count_302; // @[ToAXI4.scala 254:28]
  wire  idle_301 = ~count_302; // @[ToAXI4.scala 256:26]
  reg  count_301; // @[ToAXI4.scala 254:28]
  wire  idle_300 = ~count_301; // @[ToAXI4.scala 256:26]
  reg  count_300; // @[ToAXI4.scala 254:28]
  wire  idle_299 = ~count_300; // @[ToAXI4.scala 256:26]
  reg  count_299; // @[ToAXI4.scala 254:28]
  wire  idle_298 = ~count_299; // @[ToAXI4.scala 256:26]
  reg  count_298; // @[ToAXI4.scala 254:28]
  wire  idle_297 = ~count_298; // @[ToAXI4.scala 256:26]
  reg  count_297; // @[ToAXI4.scala 254:28]
  wire  idle_296 = ~count_297; // @[ToAXI4.scala 256:26]
  reg  count_296; // @[ToAXI4.scala 254:28]
  wire  idle_295 = ~count_296; // @[ToAXI4.scala 256:26]
  reg  count_295; // @[ToAXI4.scala 254:28]
  wire  idle_294 = ~count_295; // @[ToAXI4.scala 256:26]
  reg  count_294; // @[ToAXI4.scala 254:28]
  wire  idle_293 = ~count_294; // @[ToAXI4.scala 256:26]
  reg  count_293; // @[ToAXI4.scala 254:28]
  wire  idle_292 = ~count_293; // @[ToAXI4.scala 256:26]
  reg  count_292; // @[ToAXI4.scala 254:28]
  wire  idle_291 = ~count_292; // @[ToAXI4.scala 256:26]
  reg  count_291; // @[ToAXI4.scala 254:28]
  wire  idle_290 = ~count_291; // @[ToAXI4.scala 256:26]
  reg  count_290; // @[ToAXI4.scala 254:28]
  wire  idle_289 = ~count_290; // @[ToAXI4.scala 256:26]
  reg  count_289; // @[ToAXI4.scala 254:28]
  wire  idle_288 = ~count_289; // @[ToAXI4.scala 256:26]
  reg  count_288; // @[ToAXI4.scala 254:28]
  wire  idle_287 = ~count_288; // @[ToAXI4.scala 256:26]
  reg  count_287; // @[ToAXI4.scala 254:28]
  wire  idle_286 = ~count_287; // @[ToAXI4.scala 256:26]
  reg  count_286; // @[ToAXI4.scala 254:28]
  wire  idle_285 = ~count_286; // @[ToAXI4.scala 256:26]
  reg  count_285; // @[ToAXI4.scala 254:28]
  wire  idle_284 = ~count_285; // @[ToAXI4.scala 256:26]
  reg  count_284; // @[ToAXI4.scala 254:28]
  wire  idle_283 = ~count_284; // @[ToAXI4.scala 256:26]
  reg  count_283; // @[ToAXI4.scala 254:28]
  wire  idle_282 = ~count_283; // @[ToAXI4.scala 256:26]
  reg  count_282; // @[ToAXI4.scala 254:28]
  wire  idle_281 = ~count_282; // @[ToAXI4.scala 256:26]
  reg  count_281; // @[ToAXI4.scala 254:28]
  wire  idle_280 = ~count_281; // @[ToAXI4.scala 256:26]
  reg  count_280; // @[ToAXI4.scala 254:28]
  wire  idle_279 = ~count_280; // @[ToAXI4.scala 256:26]
  reg  count_279; // @[ToAXI4.scala 254:28]
  wire  idle_278 = ~count_279; // @[ToAXI4.scala 256:26]
  reg  count_278; // @[ToAXI4.scala 254:28]
  wire  idle_277 = ~count_278; // @[ToAXI4.scala 256:26]
  reg  count_277; // @[ToAXI4.scala 254:28]
  wire  idle_276 = ~count_277; // @[ToAXI4.scala 256:26]
  reg  count_276; // @[ToAXI4.scala 254:28]
  wire  idle_275 = ~count_276; // @[ToAXI4.scala 256:26]
  reg  count_275; // @[ToAXI4.scala 254:28]
  wire  idle_274 = ~count_275; // @[ToAXI4.scala 256:26]
  reg  count_274; // @[ToAXI4.scala 254:28]
  wire  idle_273 = ~count_274; // @[ToAXI4.scala 256:26]
  reg  count_273; // @[ToAXI4.scala 254:28]
  wire  idle_272 = ~count_273; // @[ToAXI4.scala 256:26]
  reg  count_272; // @[ToAXI4.scala 254:28]
  wire  idle_271 = ~count_272; // @[ToAXI4.scala 256:26]
  reg  count_271; // @[ToAXI4.scala 254:28]
  wire  idle_270 = ~count_271; // @[ToAXI4.scala 256:26]
  reg  count_270; // @[ToAXI4.scala 254:28]
  wire  idle_269 = ~count_270; // @[ToAXI4.scala 256:26]
  reg  count_269; // @[ToAXI4.scala 254:28]
  wire  idle_268 = ~count_269; // @[ToAXI4.scala 256:26]
  reg  count_268; // @[ToAXI4.scala 254:28]
  wire  idle_267 = ~count_268; // @[ToAXI4.scala 256:26]
  reg  count_267; // @[ToAXI4.scala 254:28]
  wire  idle_266 = ~count_267; // @[ToAXI4.scala 256:26]
  reg  count_266; // @[ToAXI4.scala 254:28]
  wire  idle_265 = ~count_266; // @[ToAXI4.scala 256:26]
  reg  count_265; // @[ToAXI4.scala 254:28]
  wire  idle_264 = ~count_265; // @[ToAXI4.scala 256:26]
  reg  count_264; // @[ToAXI4.scala 254:28]
  wire  idle_263 = ~count_264; // @[ToAXI4.scala 256:26]
  reg  count_263; // @[ToAXI4.scala 254:28]
  wire  idle_262 = ~count_263; // @[ToAXI4.scala 256:26]
  reg  count_262; // @[ToAXI4.scala 254:28]
  wire  idle_261 = ~count_262; // @[ToAXI4.scala 256:26]
  reg  count_261; // @[ToAXI4.scala 254:28]
  wire  idle_260 = ~count_261; // @[ToAXI4.scala 256:26]
  reg  count_260; // @[ToAXI4.scala 254:28]
  wire  idle_259 = ~count_260; // @[ToAXI4.scala 256:26]
  reg  count_259; // @[ToAXI4.scala 254:28]
  wire  idle_258 = ~count_259; // @[ToAXI4.scala 256:26]
  reg  count_258; // @[ToAXI4.scala 254:28]
  wire  idle_257 = ~count_258; // @[ToAXI4.scala 256:26]
  reg  count_257; // @[ToAXI4.scala 254:28]
  wire  idle_256 = ~count_257; // @[ToAXI4.scala 256:26]
  reg  count_256; // @[ToAXI4.scala 254:28]
  wire  idle_255 = ~count_256; // @[ToAXI4.scala 256:26]
  reg  count_255; // @[ToAXI4.scala 254:28]
  wire  idle_254 = ~count_255; // @[ToAXI4.scala 256:26]
  reg  count_254; // @[ToAXI4.scala 254:28]
  wire  idle_253 = ~count_254; // @[ToAXI4.scala 256:26]
  reg  count_253; // @[ToAXI4.scala 254:28]
  wire  idle_252 = ~count_253; // @[ToAXI4.scala 256:26]
  reg  count_252; // @[ToAXI4.scala 254:28]
  wire  idle_251 = ~count_252; // @[ToAXI4.scala 256:26]
  reg  count_251; // @[ToAXI4.scala 254:28]
  wire  idle_250 = ~count_251; // @[ToAXI4.scala 256:26]
  reg  count_250; // @[ToAXI4.scala 254:28]
  wire  idle_249 = ~count_250; // @[ToAXI4.scala 256:26]
  reg  count_249; // @[ToAXI4.scala 254:28]
  wire  idle_248 = ~count_249; // @[ToAXI4.scala 256:26]
  reg  count_248; // @[ToAXI4.scala 254:28]
  wire  idle_247 = ~count_248; // @[ToAXI4.scala 256:26]
  reg  count_247; // @[ToAXI4.scala 254:28]
  wire  idle_246 = ~count_247; // @[ToAXI4.scala 256:26]
  reg  count_246; // @[ToAXI4.scala 254:28]
  wire  idle_245 = ~count_246; // @[ToAXI4.scala 256:26]
  reg  count_245; // @[ToAXI4.scala 254:28]
  wire  idle_244 = ~count_245; // @[ToAXI4.scala 256:26]
  reg  count_244; // @[ToAXI4.scala 254:28]
  wire  idle_243 = ~count_244; // @[ToAXI4.scala 256:26]
  reg  count_243; // @[ToAXI4.scala 254:28]
  wire  idle_242 = ~count_243; // @[ToAXI4.scala 256:26]
  reg  count_242; // @[ToAXI4.scala 254:28]
  wire  idle_241 = ~count_242; // @[ToAXI4.scala 256:26]
  reg  count_241; // @[ToAXI4.scala 254:28]
  wire  idle_240 = ~count_241; // @[ToAXI4.scala 256:26]
  reg  count_240; // @[ToAXI4.scala 254:28]
  wire  idle_239 = ~count_240; // @[ToAXI4.scala 256:26]
  reg  count_239; // @[ToAXI4.scala 254:28]
  wire  idle_238 = ~count_239; // @[ToAXI4.scala 256:26]
  reg  count_238; // @[ToAXI4.scala 254:28]
  wire  idle_237 = ~count_238; // @[ToAXI4.scala 256:26]
  reg  count_237; // @[ToAXI4.scala 254:28]
  wire  idle_236 = ~count_237; // @[ToAXI4.scala 256:26]
  reg  count_236; // @[ToAXI4.scala 254:28]
  wire  idle_235 = ~count_236; // @[ToAXI4.scala 256:26]
  reg  count_235; // @[ToAXI4.scala 254:28]
  wire  idle_234 = ~count_235; // @[ToAXI4.scala 256:26]
  reg  count_234; // @[ToAXI4.scala 254:28]
  wire  idle_233 = ~count_234; // @[ToAXI4.scala 256:26]
  reg  count_233; // @[ToAXI4.scala 254:28]
  wire  idle_232 = ~count_233; // @[ToAXI4.scala 256:26]
  reg  count_232; // @[ToAXI4.scala 254:28]
  wire  idle_231 = ~count_232; // @[ToAXI4.scala 256:26]
  reg  count_231; // @[ToAXI4.scala 254:28]
  wire  idle_230 = ~count_231; // @[ToAXI4.scala 256:26]
  reg  count_230; // @[ToAXI4.scala 254:28]
  wire  idle_229 = ~count_230; // @[ToAXI4.scala 256:26]
  reg  count_229; // @[ToAXI4.scala 254:28]
  wire  idle_228 = ~count_229; // @[ToAXI4.scala 256:26]
  reg  count_228; // @[ToAXI4.scala 254:28]
  wire  idle_227 = ~count_228; // @[ToAXI4.scala 256:26]
  reg  count_227; // @[ToAXI4.scala 254:28]
  wire  idle_226 = ~count_227; // @[ToAXI4.scala 256:26]
  reg  count_226; // @[ToAXI4.scala 254:28]
  wire  idle_225 = ~count_226; // @[ToAXI4.scala 256:26]
  reg  count_225; // @[ToAXI4.scala 254:28]
  wire  idle_224 = ~count_225; // @[ToAXI4.scala 256:26]
  reg  count_224; // @[ToAXI4.scala 254:28]
  wire  idle_223 = ~count_224; // @[ToAXI4.scala 256:26]
  reg  count_223; // @[ToAXI4.scala 254:28]
  wire  idle_222 = ~count_223; // @[ToAXI4.scala 256:26]
  reg  count_222; // @[ToAXI4.scala 254:28]
  wire  idle_221 = ~count_222; // @[ToAXI4.scala 256:26]
  reg  count_221; // @[ToAXI4.scala 254:28]
  wire  idle_220 = ~count_221; // @[ToAXI4.scala 256:26]
  reg  count_220; // @[ToAXI4.scala 254:28]
  wire  idle_219 = ~count_220; // @[ToAXI4.scala 256:26]
  reg  count_219; // @[ToAXI4.scala 254:28]
  wire  idle_218 = ~count_219; // @[ToAXI4.scala 256:26]
  reg  count_218; // @[ToAXI4.scala 254:28]
  wire  idle_217 = ~count_218; // @[ToAXI4.scala 256:26]
  reg  count_217; // @[ToAXI4.scala 254:28]
  wire  idle_216 = ~count_217; // @[ToAXI4.scala 256:26]
  reg  count_216; // @[ToAXI4.scala 254:28]
  wire  idle_215 = ~count_216; // @[ToAXI4.scala 256:26]
  reg  count_215; // @[ToAXI4.scala 254:28]
  wire  idle_214 = ~count_215; // @[ToAXI4.scala 256:26]
  reg  count_214; // @[ToAXI4.scala 254:28]
  wire  idle_213 = ~count_214; // @[ToAXI4.scala 256:26]
  reg  count_213; // @[ToAXI4.scala 254:28]
  wire  idle_212 = ~count_213; // @[ToAXI4.scala 256:26]
  reg  count_212; // @[ToAXI4.scala 254:28]
  wire  idle_211 = ~count_212; // @[ToAXI4.scala 256:26]
  reg  count_211; // @[ToAXI4.scala 254:28]
  wire  idle_210 = ~count_211; // @[ToAXI4.scala 256:26]
  reg  count_210; // @[ToAXI4.scala 254:28]
  wire  idle_209 = ~count_210; // @[ToAXI4.scala 256:26]
  reg  count_209; // @[ToAXI4.scala 254:28]
  wire  idle_208 = ~count_209; // @[ToAXI4.scala 256:26]
  reg  count_208; // @[ToAXI4.scala 254:28]
  wire  idle_207 = ~count_208; // @[ToAXI4.scala 256:26]
  reg  count_207; // @[ToAXI4.scala 254:28]
  wire  idle_206 = ~count_207; // @[ToAXI4.scala 256:26]
  reg  count_206; // @[ToAXI4.scala 254:28]
  wire  idle_205 = ~count_206; // @[ToAXI4.scala 256:26]
  reg  count_205; // @[ToAXI4.scala 254:28]
  wire  idle_204 = ~count_205; // @[ToAXI4.scala 256:26]
  reg  count_204; // @[ToAXI4.scala 254:28]
  wire  idle_203 = ~count_204; // @[ToAXI4.scala 256:26]
  reg  count_203; // @[ToAXI4.scala 254:28]
  wire  idle_202 = ~count_203; // @[ToAXI4.scala 256:26]
  reg  count_202; // @[ToAXI4.scala 254:28]
  wire  idle_201 = ~count_202; // @[ToAXI4.scala 256:26]
  reg  count_201; // @[ToAXI4.scala 254:28]
  wire  idle_200 = ~count_201; // @[ToAXI4.scala 256:26]
  reg  count_200; // @[ToAXI4.scala 254:28]
  wire  idle_199 = ~count_200; // @[ToAXI4.scala 256:26]
  reg  count_199; // @[ToAXI4.scala 254:28]
  wire  idle_198 = ~count_199; // @[ToAXI4.scala 256:26]
  reg  count_198; // @[ToAXI4.scala 254:28]
  wire  idle_197 = ~count_198; // @[ToAXI4.scala 256:26]
  reg  count_197; // @[ToAXI4.scala 254:28]
  wire  idle_196 = ~count_197; // @[ToAXI4.scala 256:26]
  reg  count_196; // @[ToAXI4.scala 254:28]
  wire  idle_195 = ~count_196; // @[ToAXI4.scala 256:26]
  reg  count_195; // @[ToAXI4.scala 254:28]
  wire  idle_194 = ~count_195; // @[ToAXI4.scala 256:26]
  reg  count_194; // @[ToAXI4.scala 254:28]
  wire  idle_193 = ~count_194; // @[ToAXI4.scala 256:26]
  reg  count_193; // @[ToAXI4.scala 254:28]
  wire  idle_192 = ~count_193; // @[ToAXI4.scala 256:26]
  reg  count_192; // @[ToAXI4.scala 254:28]
  wire  idle_191 = ~count_192; // @[ToAXI4.scala 256:26]
  reg  count_191; // @[ToAXI4.scala 254:28]
  wire  idle_190 = ~count_191; // @[ToAXI4.scala 256:26]
  reg  count_190; // @[ToAXI4.scala 254:28]
  wire  idle_189 = ~count_190; // @[ToAXI4.scala 256:26]
  reg  count_189; // @[ToAXI4.scala 254:28]
  wire  idle_188 = ~count_189; // @[ToAXI4.scala 256:26]
  reg  count_188; // @[ToAXI4.scala 254:28]
  wire  idle_187 = ~count_188; // @[ToAXI4.scala 256:26]
  reg  count_187; // @[ToAXI4.scala 254:28]
  wire  idle_186 = ~count_187; // @[ToAXI4.scala 256:26]
  reg  count_186; // @[ToAXI4.scala 254:28]
  wire  idle_185 = ~count_186; // @[ToAXI4.scala 256:26]
  reg  count_185; // @[ToAXI4.scala 254:28]
  wire  idle_184 = ~count_185; // @[ToAXI4.scala 256:26]
  reg  count_184; // @[ToAXI4.scala 254:28]
  wire  idle_183 = ~count_184; // @[ToAXI4.scala 256:26]
  reg  count_183; // @[ToAXI4.scala 254:28]
  wire  idle_182 = ~count_183; // @[ToAXI4.scala 256:26]
  reg  count_182; // @[ToAXI4.scala 254:28]
  wire  idle_181 = ~count_182; // @[ToAXI4.scala 256:26]
  reg  count_181; // @[ToAXI4.scala 254:28]
  wire  idle_180 = ~count_181; // @[ToAXI4.scala 256:26]
  reg  count_180; // @[ToAXI4.scala 254:28]
  wire  idle_179 = ~count_180; // @[ToAXI4.scala 256:26]
  reg  count_179; // @[ToAXI4.scala 254:28]
  wire  idle_178 = ~count_179; // @[ToAXI4.scala 256:26]
  reg  count_178; // @[ToAXI4.scala 254:28]
  wire  idle_177 = ~count_178; // @[ToAXI4.scala 256:26]
  reg  count_177; // @[ToAXI4.scala 254:28]
  wire  idle_176 = ~count_177; // @[ToAXI4.scala 256:26]
  reg  count_176; // @[ToAXI4.scala 254:28]
  wire  idle_175 = ~count_176; // @[ToAXI4.scala 256:26]
  reg  count_175; // @[ToAXI4.scala 254:28]
  wire  idle_174 = ~count_175; // @[ToAXI4.scala 256:26]
  reg  count_174; // @[ToAXI4.scala 254:28]
  wire  idle_173 = ~count_174; // @[ToAXI4.scala 256:26]
  reg  count_173; // @[ToAXI4.scala 254:28]
  wire  idle_172 = ~count_173; // @[ToAXI4.scala 256:26]
  reg  count_172; // @[ToAXI4.scala 254:28]
  wire  idle_171 = ~count_172; // @[ToAXI4.scala 256:26]
  reg  count_171; // @[ToAXI4.scala 254:28]
  wire  idle_170 = ~count_171; // @[ToAXI4.scala 256:26]
  reg  count_170; // @[ToAXI4.scala 254:28]
  wire  idle_169 = ~count_170; // @[ToAXI4.scala 256:26]
  reg  count_169; // @[ToAXI4.scala 254:28]
  wire  idle_168 = ~count_169; // @[ToAXI4.scala 256:26]
  reg  count_168; // @[ToAXI4.scala 254:28]
  wire  idle_167 = ~count_168; // @[ToAXI4.scala 256:26]
  reg  count_167; // @[ToAXI4.scala 254:28]
  wire  idle_166 = ~count_167; // @[ToAXI4.scala 256:26]
  reg  count_166; // @[ToAXI4.scala 254:28]
  wire  idle_165 = ~count_166; // @[ToAXI4.scala 256:26]
  reg  count_165; // @[ToAXI4.scala 254:28]
  wire  idle_164 = ~count_165; // @[ToAXI4.scala 256:26]
  reg  count_164; // @[ToAXI4.scala 254:28]
  wire  idle_163 = ~count_164; // @[ToAXI4.scala 256:26]
  reg  count_163; // @[ToAXI4.scala 254:28]
  wire  idle_162 = ~count_163; // @[ToAXI4.scala 256:26]
  reg  count_162; // @[ToAXI4.scala 254:28]
  wire  idle_161 = ~count_162; // @[ToAXI4.scala 256:26]
  reg  count_161; // @[ToAXI4.scala 254:28]
  wire  idle_160 = ~count_161; // @[ToAXI4.scala 256:26]
  reg  count_160; // @[ToAXI4.scala 254:28]
  wire  idle_159 = ~count_160; // @[ToAXI4.scala 256:26]
  reg  count_159; // @[ToAXI4.scala 254:28]
  wire  idle_158 = ~count_159; // @[ToAXI4.scala 256:26]
  reg  count_158; // @[ToAXI4.scala 254:28]
  wire  idle_157 = ~count_158; // @[ToAXI4.scala 256:26]
  reg  count_157; // @[ToAXI4.scala 254:28]
  wire  idle_156 = ~count_157; // @[ToAXI4.scala 256:26]
  reg  count_156; // @[ToAXI4.scala 254:28]
  wire  idle_155 = ~count_156; // @[ToAXI4.scala 256:26]
  reg  count_155; // @[ToAXI4.scala 254:28]
  wire  idle_154 = ~count_155; // @[ToAXI4.scala 256:26]
  reg  count_154; // @[ToAXI4.scala 254:28]
  wire  idle_153 = ~count_154; // @[ToAXI4.scala 256:26]
  reg  count_153; // @[ToAXI4.scala 254:28]
  wire  idle_152 = ~count_153; // @[ToAXI4.scala 256:26]
  reg  count_152; // @[ToAXI4.scala 254:28]
  wire  idle_151 = ~count_152; // @[ToAXI4.scala 256:26]
  reg  count_151; // @[ToAXI4.scala 254:28]
  wire  idle_150 = ~count_151; // @[ToAXI4.scala 256:26]
  reg  count_150; // @[ToAXI4.scala 254:28]
  wire  idle_149 = ~count_150; // @[ToAXI4.scala 256:26]
  reg  count_149; // @[ToAXI4.scala 254:28]
  wire  idle_148 = ~count_149; // @[ToAXI4.scala 256:26]
  reg  count_148; // @[ToAXI4.scala 254:28]
  wire  idle_147 = ~count_148; // @[ToAXI4.scala 256:26]
  reg  count_147; // @[ToAXI4.scala 254:28]
  wire  idle_146 = ~count_147; // @[ToAXI4.scala 256:26]
  reg  count_146; // @[ToAXI4.scala 254:28]
  wire  idle_145 = ~count_146; // @[ToAXI4.scala 256:26]
  reg  count_145; // @[ToAXI4.scala 254:28]
  wire  idle_144 = ~count_145; // @[ToAXI4.scala 256:26]
  reg  count_144; // @[ToAXI4.scala 254:28]
  wire  idle_143 = ~count_144; // @[ToAXI4.scala 256:26]
  reg  count_143; // @[ToAXI4.scala 254:28]
  wire  idle_142 = ~count_143; // @[ToAXI4.scala 256:26]
  reg  count_142; // @[ToAXI4.scala 254:28]
  wire  idle_141 = ~count_142; // @[ToAXI4.scala 256:26]
  reg  count_141; // @[ToAXI4.scala 254:28]
  wire  idle_140 = ~count_141; // @[ToAXI4.scala 256:26]
  reg  count_140; // @[ToAXI4.scala 254:28]
  wire  idle_139 = ~count_140; // @[ToAXI4.scala 256:26]
  reg  count_139; // @[ToAXI4.scala 254:28]
  wire  idle_138 = ~count_139; // @[ToAXI4.scala 256:26]
  reg  count_138; // @[ToAXI4.scala 254:28]
  wire  idle_137 = ~count_138; // @[ToAXI4.scala 256:26]
  reg  count_137; // @[ToAXI4.scala 254:28]
  wire  idle_136 = ~count_137; // @[ToAXI4.scala 256:26]
  reg  count_136; // @[ToAXI4.scala 254:28]
  wire  idle_135 = ~count_136; // @[ToAXI4.scala 256:26]
  reg  count_135; // @[ToAXI4.scala 254:28]
  wire  idle_134 = ~count_135; // @[ToAXI4.scala 256:26]
  reg  count_134; // @[ToAXI4.scala 254:28]
  wire  idle_133 = ~count_134; // @[ToAXI4.scala 256:26]
  reg  count_133; // @[ToAXI4.scala 254:28]
  wire  idle_132 = ~count_133; // @[ToAXI4.scala 256:26]
  reg  count_132; // @[ToAXI4.scala 254:28]
  wire  idle_131 = ~count_132; // @[ToAXI4.scala 256:26]
  reg  count_131; // @[ToAXI4.scala 254:28]
  wire  idle_130 = ~count_131; // @[ToAXI4.scala 256:26]
  reg  count_130; // @[ToAXI4.scala 254:28]
  wire  idle_129 = ~count_130; // @[ToAXI4.scala 256:26]
  reg  count_129; // @[ToAXI4.scala 254:28]
  wire  idle_128 = ~count_129; // @[ToAXI4.scala 256:26]
  reg  count_128; // @[ToAXI4.scala 254:28]
  wire  idle_127 = ~count_128; // @[ToAXI4.scala 256:26]
  reg  count_127; // @[ToAXI4.scala 254:28]
  wire  idle_126 = ~count_127; // @[ToAXI4.scala 256:26]
  reg  count_126; // @[ToAXI4.scala 254:28]
  wire  idle_125 = ~count_126; // @[ToAXI4.scala 256:26]
  reg  count_125; // @[ToAXI4.scala 254:28]
  wire  idle_124 = ~count_125; // @[ToAXI4.scala 256:26]
  reg  count_124; // @[ToAXI4.scala 254:28]
  wire  idle_123 = ~count_124; // @[ToAXI4.scala 256:26]
  reg  count_123; // @[ToAXI4.scala 254:28]
  wire  idle_122 = ~count_123; // @[ToAXI4.scala 256:26]
  reg  count_122; // @[ToAXI4.scala 254:28]
  wire  idle_121 = ~count_122; // @[ToAXI4.scala 256:26]
  reg  count_121; // @[ToAXI4.scala 254:28]
  wire  idle_120 = ~count_121; // @[ToAXI4.scala 256:26]
  reg  count_120; // @[ToAXI4.scala 254:28]
  wire  idle_119 = ~count_120; // @[ToAXI4.scala 256:26]
  reg  count_119; // @[ToAXI4.scala 254:28]
  wire  idle_118 = ~count_119; // @[ToAXI4.scala 256:26]
  reg  count_118; // @[ToAXI4.scala 254:28]
  wire  idle_117 = ~count_118; // @[ToAXI4.scala 256:26]
  reg  count_117; // @[ToAXI4.scala 254:28]
  wire  idle_116 = ~count_117; // @[ToAXI4.scala 256:26]
  reg  count_116; // @[ToAXI4.scala 254:28]
  wire  idle_115 = ~count_116; // @[ToAXI4.scala 256:26]
  reg  count_115; // @[ToAXI4.scala 254:28]
  wire  idle_114 = ~count_115; // @[ToAXI4.scala 256:26]
  reg  count_114; // @[ToAXI4.scala 254:28]
  wire  idle_113 = ~count_114; // @[ToAXI4.scala 256:26]
  reg  count_113; // @[ToAXI4.scala 254:28]
  wire  idle_112 = ~count_113; // @[ToAXI4.scala 256:26]
  reg  count_112; // @[ToAXI4.scala 254:28]
  wire  idle_111 = ~count_112; // @[ToAXI4.scala 256:26]
  reg  count_111; // @[ToAXI4.scala 254:28]
  wire  idle_110 = ~count_111; // @[ToAXI4.scala 256:26]
  reg  count_110; // @[ToAXI4.scala 254:28]
  wire  idle_109 = ~count_110; // @[ToAXI4.scala 256:26]
  reg  count_109; // @[ToAXI4.scala 254:28]
  wire  idle_108 = ~count_109; // @[ToAXI4.scala 256:26]
  reg  count_108; // @[ToAXI4.scala 254:28]
  wire  idle_107 = ~count_108; // @[ToAXI4.scala 256:26]
  reg  count_107; // @[ToAXI4.scala 254:28]
  wire  idle_106 = ~count_107; // @[ToAXI4.scala 256:26]
  reg  count_106; // @[ToAXI4.scala 254:28]
  wire  idle_105 = ~count_106; // @[ToAXI4.scala 256:26]
  reg  count_105; // @[ToAXI4.scala 254:28]
  wire  idle_104 = ~count_105; // @[ToAXI4.scala 256:26]
  reg  count_104; // @[ToAXI4.scala 254:28]
  wire  idle_103 = ~count_104; // @[ToAXI4.scala 256:26]
  reg  count_103; // @[ToAXI4.scala 254:28]
  wire  idle_102 = ~count_103; // @[ToAXI4.scala 256:26]
  reg  count_102; // @[ToAXI4.scala 254:28]
  wire  idle_101 = ~count_102; // @[ToAXI4.scala 256:26]
  reg  count_101; // @[ToAXI4.scala 254:28]
  wire  idle_100 = ~count_101; // @[ToAXI4.scala 256:26]
  reg  count_100; // @[ToAXI4.scala 254:28]
  wire  idle_99 = ~count_100; // @[ToAXI4.scala 256:26]
  reg  count_99; // @[ToAXI4.scala 254:28]
  wire  idle_98 = ~count_99; // @[ToAXI4.scala 256:26]
  reg  count_98; // @[ToAXI4.scala 254:28]
  wire  idle_97 = ~count_98; // @[ToAXI4.scala 256:26]
  reg  count_97; // @[ToAXI4.scala 254:28]
  wire  idle_96 = ~count_97; // @[ToAXI4.scala 256:26]
  reg  count_96; // @[ToAXI4.scala 254:28]
  wire  idle_95 = ~count_96; // @[ToAXI4.scala 256:26]
  reg  count_95; // @[ToAXI4.scala 254:28]
  wire  idle_94 = ~count_95; // @[ToAXI4.scala 256:26]
  reg  count_94; // @[ToAXI4.scala 254:28]
  wire  idle_93 = ~count_94; // @[ToAXI4.scala 256:26]
  reg  count_93; // @[ToAXI4.scala 254:28]
  wire  idle_92 = ~count_93; // @[ToAXI4.scala 256:26]
  reg  count_92; // @[ToAXI4.scala 254:28]
  wire  idle_91 = ~count_92; // @[ToAXI4.scala 256:26]
  reg  count_91; // @[ToAXI4.scala 254:28]
  wire  idle_90 = ~count_91; // @[ToAXI4.scala 256:26]
  reg  count_90; // @[ToAXI4.scala 254:28]
  wire  idle_89 = ~count_90; // @[ToAXI4.scala 256:26]
  reg  count_89; // @[ToAXI4.scala 254:28]
  wire  idle_88 = ~count_89; // @[ToAXI4.scala 256:26]
  reg  count_88; // @[ToAXI4.scala 254:28]
  wire  idle_87 = ~count_88; // @[ToAXI4.scala 256:26]
  reg  count_87; // @[ToAXI4.scala 254:28]
  wire  idle_86 = ~count_87; // @[ToAXI4.scala 256:26]
  reg  count_86; // @[ToAXI4.scala 254:28]
  wire  idle_85 = ~count_86; // @[ToAXI4.scala 256:26]
  reg  count_85; // @[ToAXI4.scala 254:28]
  wire  idle_84 = ~count_85; // @[ToAXI4.scala 256:26]
  reg  count_84; // @[ToAXI4.scala 254:28]
  wire  idle_83 = ~count_84; // @[ToAXI4.scala 256:26]
  reg  count_83; // @[ToAXI4.scala 254:28]
  wire  idle_82 = ~count_83; // @[ToAXI4.scala 256:26]
  reg  count_82; // @[ToAXI4.scala 254:28]
  wire  idle_81 = ~count_82; // @[ToAXI4.scala 256:26]
  reg  count_81; // @[ToAXI4.scala 254:28]
  wire  idle_80 = ~count_81; // @[ToAXI4.scala 256:26]
  reg  count_80; // @[ToAXI4.scala 254:28]
  wire  idle_79 = ~count_80; // @[ToAXI4.scala 256:26]
  reg  count_79; // @[ToAXI4.scala 254:28]
  wire  idle_78 = ~count_79; // @[ToAXI4.scala 256:26]
  reg  count_78; // @[ToAXI4.scala 254:28]
  wire  idle_77 = ~count_78; // @[ToAXI4.scala 256:26]
  reg  count_77; // @[ToAXI4.scala 254:28]
  wire  idle_76 = ~count_77; // @[ToAXI4.scala 256:26]
  reg  count_76; // @[ToAXI4.scala 254:28]
  wire  idle_75 = ~count_76; // @[ToAXI4.scala 256:26]
  reg  count_75; // @[ToAXI4.scala 254:28]
  wire  idle_74 = ~count_75; // @[ToAXI4.scala 256:26]
  reg  count_74; // @[ToAXI4.scala 254:28]
  wire  idle_73 = ~count_74; // @[ToAXI4.scala 256:26]
  reg  count_73; // @[ToAXI4.scala 254:28]
  wire  idle_72 = ~count_73; // @[ToAXI4.scala 256:26]
  reg  count_72; // @[ToAXI4.scala 254:28]
  wire  idle_71 = ~count_72; // @[ToAXI4.scala 256:26]
  reg  count_71; // @[ToAXI4.scala 254:28]
  wire  idle_70 = ~count_71; // @[ToAXI4.scala 256:26]
  reg  count_70; // @[ToAXI4.scala 254:28]
  wire  idle_69 = ~count_70; // @[ToAXI4.scala 256:26]
  reg  count_69; // @[ToAXI4.scala 254:28]
  wire  idle_68 = ~count_69; // @[ToAXI4.scala 256:26]
  reg  count_68; // @[ToAXI4.scala 254:28]
  wire  idle_67 = ~count_68; // @[ToAXI4.scala 256:26]
  reg  count_67; // @[ToAXI4.scala 254:28]
  wire  idle_66 = ~count_67; // @[ToAXI4.scala 256:26]
  reg  count_66; // @[ToAXI4.scala 254:28]
  wire  idle_65 = ~count_66; // @[ToAXI4.scala 256:26]
  reg  count_65; // @[ToAXI4.scala 254:28]
  wire  idle_64 = ~count_65; // @[ToAXI4.scala 256:26]
  reg  count_64; // @[ToAXI4.scala 254:28]
  wire  idle_63 = ~count_64; // @[ToAXI4.scala 256:26]
  reg  count_63; // @[ToAXI4.scala 254:28]
  wire  idle_62 = ~count_63; // @[ToAXI4.scala 256:26]
  reg  count_62; // @[ToAXI4.scala 254:28]
  wire  idle_61 = ~count_62; // @[ToAXI4.scala 256:26]
  reg  count_61; // @[ToAXI4.scala 254:28]
  wire  idle_60 = ~count_61; // @[ToAXI4.scala 256:26]
  reg  count_60; // @[ToAXI4.scala 254:28]
  wire  idle_59 = ~count_60; // @[ToAXI4.scala 256:26]
  reg  count_59; // @[ToAXI4.scala 254:28]
  wire  idle_58 = ~count_59; // @[ToAXI4.scala 256:26]
  reg  count_58; // @[ToAXI4.scala 254:28]
  wire  idle_57 = ~count_58; // @[ToAXI4.scala 256:26]
  reg  count_57; // @[ToAXI4.scala 254:28]
  wire  idle_56 = ~count_57; // @[ToAXI4.scala 256:26]
  reg  count_56; // @[ToAXI4.scala 254:28]
  wire  idle_55 = ~count_56; // @[ToAXI4.scala 256:26]
  reg  count_55; // @[ToAXI4.scala 254:28]
  wire  idle_54 = ~count_55; // @[ToAXI4.scala 256:26]
  reg  count_54; // @[ToAXI4.scala 254:28]
  wire  idle_53 = ~count_54; // @[ToAXI4.scala 256:26]
  reg  count_53; // @[ToAXI4.scala 254:28]
  wire  idle_52 = ~count_53; // @[ToAXI4.scala 256:26]
  reg  count_52; // @[ToAXI4.scala 254:28]
  wire  idle_51 = ~count_52; // @[ToAXI4.scala 256:26]
  reg  count_51; // @[ToAXI4.scala 254:28]
  wire  idle_50 = ~count_51; // @[ToAXI4.scala 256:26]
  reg  count_50; // @[ToAXI4.scala 254:28]
  wire  idle_49 = ~count_50; // @[ToAXI4.scala 256:26]
  reg  count_49; // @[ToAXI4.scala 254:28]
  wire  idle_48 = ~count_49; // @[ToAXI4.scala 256:26]
  reg  count_48; // @[ToAXI4.scala 254:28]
  wire  idle_47 = ~count_48; // @[ToAXI4.scala 256:26]
  reg  count_47; // @[ToAXI4.scala 254:28]
  wire  idle_46 = ~count_47; // @[ToAXI4.scala 256:26]
  reg  count_46; // @[ToAXI4.scala 254:28]
  wire  idle_45 = ~count_46; // @[ToAXI4.scala 256:26]
  reg  count_45; // @[ToAXI4.scala 254:28]
  wire  idle_44 = ~count_45; // @[ToAXI4.scala 256:26]
  reg  count_44; // @[ToAXI4.scala 254:28]
  wire  idle_43 = ~count_44; // @[ToAXI4.scala 256:26]
  reg  count_43; // @[ToAXI4.scala 254:28]
  wire  idle_42 = ~count_43; // @[ToAXI4.scala 256:26]
  reg  count_42; // @[ToAXI4.scala 254:28]
  wire  idle_41 = ~count_42; // @[ToAXI4.scala 256:26]
  reg  count_41; // @[ToAXI4.scala 254:28]
  wire  idle_40 = ~count_41; // @[ToAXI4.scala 256:26]
  reg  count_40; // @[ToAXI4.scala 254:28]
  wire  idle_39 = ~count_40; // @[ToAXI4.scala 256:26]
  reg  count_39; // @[ToAXI4.scala 254:28]
  wire  idle_38 = ~count_39; // @[ToAXI4.scala 256:26]
  reg  count_38; // @[ToAXI4.scala 254:28]
  wire  idle_37 = ~count_38; // @[ToAXI4.scala 256:26]
  reg  count_37; // @[ToAXI4.scala 254:28]
  wire  idle_36 = ~count_37; // @[ToAXI4.scala 256:26]
  reg  count_36; // @[ToAXI4.scala 254:28]
  wire  idle_35 = ~count_36; // @[ToAXI4.scala 256:26]
  reg  count_35; // @[ToAXI4.scala 254:28]
  wire  idle_34 = ~count_35; // @[ToAXI4.scala 256:26]
  reg  count_34; // @[ToAXI4.scala 254:28]
  wire  idle_33 = ~count_34; // @[ToAXI4.scala 256:26]
  reg  count_33; // @[ToAXI4.scala 254:28]
  wire  idle_32 = ~count_33; // @[ToAXI4.scala 256:26]
  reg  count_32; // @[ToAXI4.scala 254:28]
  wire  idle_31 = ~count_32; // @[ToAXI4.scala 256:26]
  reg  count_31; // @[ToAXI4.scala 254:28]
  wire  idle_30 = ~count_31; // @[ToAXI4.scala 256:26]
  reg  count_30; // @[ToAXI4.scala 254:28]
  wire  idle_29 = ~count_30; // @[ToAXI4.scala 256:26]
  reg  count_29; // @[ToAXI4.scala 254:28]
  wire  idle_28 = ~count_29; // @[ToAXI4.scala 256:26]
  reg  count_28; // @[ToAXI4.scala 254:28]
  wire  idle_27 = ~count_28; // @[ToAXI4.scala 256:26]
  reg  count_27; // @[ToAXI4.scala 254:28]
  wire  idle_26 = ~count_27; // @[ToAXI4.scala 256:26]
  reg  count_26; // @[ToAXI4.scala 254:28]
  wire  idle_25 = ~count_26; // @[ToAXI4.scala 256:26]
  reg  count_25; // @[ToAXI4.scala 254:28]
  wire  idle_24 = ~count_25; // @[ToAXI4.scala 256:26]
  reg  count_24; // @[ToAXI4.scala 254:28]
  wire  idle_23 = ~count_24; // @[ToAXI4.scala 256:26]
  reg  count_23; // @[ToAXI4.scala 254:28]
  wire  idle_22 = ~count_23; // @[ToAXI4.scala 256:26]
  reg  count_22; // @[ToAXI4.scala 254:28]
  wire  idle_21 = ~count_22; // @[ToAXI4.scala 256:26]
  reg  count_21; // @[ToAXI4.scala 254:28]
  wire  idle_20 = ~count_21; // @[ToAXI4.scala 256:26]
  reg  count_20; // @[ToAXI4.scala 254:28]
  wire  idle_19 = ~count_20; // @[ToAXI4.scala 256:26]
  reg  count_19; // @[ToAXI4.scala 254:28]
  wire  idle_18 = ~count_19; // @[ToAXI4.scala 256:26]
  reg  count_18; // @[ToAXI4.scala 254:28]
  wire  idle_17 = ~count_18; // @[ToAXI4.scala 256:26]
  reg  count_17; // @[ToAXI4.scala 254:28]
  wire  idle_16 = ~count_17; // @[ToAXI4.scala 256:26]
  reg  count_16; // @[ToAXI4.scala 254:28]
  wire  idle_15 = ~count_16; // @[ToAXI4.scala 256:26]
  reg  count_15; // @[ToAXI4.scala 254:28]
  wire  idle_14 = ~count_15; // @[ToAXI4.scala 256:26]
  reg  count_14; // @[ToAXI4.scala 254:28]
  wire  idle_13 = ~count_14; // @[ToAXI4.scala 256:26]
  reg  count_13; // @[ToAXI4.scala 254:28]
  wire  idle_12 = ~count_13; // @[ToAXI4.scala 256:26]
  reg  count_12; // @[ToAXI4.scala 254:28]
  wire  idle_11 = ~count_12; // @[ToAXI4.scala 256:26]
  reg  count_11; // @[ToAXI4.scala 254:28]
  wire  idle_10 = ~count_11; // @[ToAXI4.scala 256:26]
  reg  count_10; // @[ToAXI4.scala 254:28]
  wire  idle_9 = ~count_10; // @[ToAXI4.scala 256:26]
  reg  count_9; // @[ToAXI4.scala 254:28]
  wire  idle_8 = ~count_9; // @[ToAXI4.scala 256:26]
  reg  count_8; // @[ToAXI4.scala 254:28]
  wire  idle_7 = ~count_8; // @[ToAXI4.scala 256:26]
  reg  count_7; // @[ToAXI4.scala 254:28]
  wire  idle_6 = ~count_7; // @[ToAXI4.scala 256:26]
  reg  count_6; // @[ToAXI4.scala 254:28]
  wire  idle_5 = ~count_6; // @[ToAXI4.scala 256:26]
  reg  count_5; // @[ToAXI4.scala 254:28]
  wire  idle_4 = ~count_5; // @[ToAXI4.scala 256:26]
  reg  count_4; // @[ToAXI4.scala 254:28]
  wire  idle_3 = ~count_4; // @[ToAXI4.scala 256:26]
  reg  count_3; // @[ToAXI4.scala 254:28]
  wire  idle_2 = ~count_3; // @[ToAXI4.scala 256:26]
  reg  count_2; // @[ToAXI4.scala 254:28]
  wire  idle_1 = ~count_2; // @[ToAXI4.scala 256:26]
  reg  count_1; // @[ToAXI4.scala 254:28]
  wire  idle = ~count_1; // @[ToAXI4.scala 256:26]
  wire  _GEN_515 = 9'h1 == auto_in_a_bits_source ? count_2 : count_1; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_516 = 9'h2 == auto_in_a_bits_source ? count_3 : _GEN_515; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_517 = 9'h3 == auto_in_a_bits_source ? count_4 : _GEN_516; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_518 = 9'h4 == auto_in_a_bits_source ? count_5 : _GEN_517; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_519 = 9'h5 == auto_in_a_bits_source ? count_6 : _GEN_518; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_520 = 9'h6 == auto_in_a_bits_source ? count_7 : _GEN_519; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_521 = 9'h7 == auto_in_a_bits_source ? count_8 : _GEN_520; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_522 = 9'h8 == auto_in_a_bits_source ? count_9 : _GEN_521; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_523 = 9'h9 == auto_in_a_bits_source ? count_10 : _GEN_522; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_524 = 9'ha == auto_in_a_bits_source ? count_11 : _GEN_523; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_525 = 9'hb == auto_in_a_bits_source ? count_12 : _GEN_524; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_526 = 9'hc == auto_in_a_bits_source ? count_13 : _GEN_525; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_527 = 9'hd == auto_in_a_bits_source ? count_14 : _GEN_526; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_528 = 9'he == auto_in_a_bits_source ? count_15 : _GEN_527; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_529 = 9'hf == auto_in_a_bits_source ? count_16 : _GEN_528; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_530 = 9'h10 == auto_in_a_bits_source ? count_17 : _GEN_529; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_531 = 9'h11 == auto_in_a_bits_source ? count_18 : _GEN_530; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_532 = 9'h12 == auto_in_a_bits_source ? count_19 : _GEN_531; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_533 = 9'h13 == auto_in_a_bits_source ? count_20 : _GEN_532; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_534 = 9'h14 == auto_in_a_bits_source ? count_21 : _GEN_533; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_535 = 9'h15 == auto_in_a_bits_source ? count_22 : _GEN_534; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_536 = 9'h16 == auto_in_a_bits_source ? count_23 : _GEN_535; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_537 = 9'h17 == auto_in_a_bits_source ? count_24 : _GEN_536; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_538 = 9'h18 == auto_in_a_bits_source ? count_25 : _GEN_537; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_539 = 9'h19 == auto_in_a_bits_source ? count_26 : _GEN_538; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_540 = 9'h1a == auto_in_a_bits_source ? count_27 : _GEN_539; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_541 = 9'h1b == auto_in_a_bits_source ? count_28 : _GEN_540; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_542 = 9'h1c == auto_in_a_bits_source ? count_29 : _GEN_541; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_543 = 9'h1d == auto_in_a_bits_source ? count_30 : _GEN_542; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_544 = 9'h1e == auto_in_a_bits_source ? count_31 : _GEN_543; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_545 = 9'h1f == auto_in_a_bits_source ? count_32 : _GEN_544; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_546 = 9'h20 == auto_in_a_bits_source ? count_33 : _GEN_545; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_547 = 9'h21 == auto_in_a_bits_source ? count_34 : _GEN_546; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_548 = 9'h22 == auto_in_a_bits_source ? count_35 : _GEN_547; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_549 = 9'h23 == auto_in_a_bits_source ? count_36 : _GEN_548; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_550 = 9'h24 == auto_in_a_bits_source ? count_37 : _GEN_549; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_551 = 9'h25 == auto_in_a_bits_source ? count_38 : _GEN_550; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_552 = 9'h26 == auto_in_a_bits_source ? count_39 : _GEN_551; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_553 = 9'h27 == auto_in_a_bits_source ? count_40 : _GEN_552; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_554 = 9'h28 == auto_in_a_bits_source ? count_41 : _GEN_553; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_555 = 9'h29 == auto_in_a_bits_source ? count_42 : _GEN_554; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_556 = 9'h2a == auto_in_a_bits_source ? count_43 : _GEN_555; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_557 = 9'h2b == auto_in_a_bits_source ? count_44 : _GEN_556; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_558 = 9'h2c == auto_in_a_bits_source ? count_45 : _GEN_557; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_559 = 9'h2d == auto_in_a_bits_source ? count_46 : _GEN_558; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_560 = 9'h2e == auto_in_a_bits_source ? count_47 : _GEN_559; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_561 = 9'h2f == auto_in_a_bits_source ? count_48 : _GEN_560; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_562 = 9'h30 == auto_in_a_bits_source ? count_49 : _GEN_561; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_563 = 9'h31 == auto_in_a_bits_source ? count_50 : _GEN_562; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_564 = 9'h32 == auto_in_a_bits_source ? count_51 : _GEN_563; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_565 = 9'h33 == auto_in_a_bits_source ? count_52 : _GEN_564; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_566 = 9'h34 == auto_in_a_bits_source ? count_53 : _GEN_565; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_567 = 9'h35 == auto_in_a_bits_source ? count_54 : _GEN_566; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_568 = 9'h36 == auto_in_a_bits_source ? count_55 : _GEN_567; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_569 = 9'h37 == auto_in_a_bits_source ? count_56 : _GEN_568; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_570 = 9'h38 == auto_in_a_bits_source ? count_57 : _GEN_569; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_571 = 9'h39 == auto_in_a_bits_source ? count_58 : _GEN_570; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_572 = 9'h3a == auto_in_a_bits_source ? count_59 : _GEN_571; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_573 = 9'h3b == auto_in_a_bits_source ? count_60 : _GEN_572; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_574 = 9'h3c == auto_in_a_bits_source ? count_61 : _GEN_573; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_575 = 9'h3d == auto_in_a_bits_source ? count_62 : _GEN_574; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_576 = 9'h3e == auto_in_a_bits_source ? count_63 : _GEN_575; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_577 = 9'h3f == auto_in_a_bits_source ? count_64 : _GEN_576; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_578 = 9'h40 == auto_in_a_bits_source ? count_65 : _GEN_577; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_579 = 9'h41 == auto_in_a_bits_source ? count_66 : _GEN_578; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_580 = 9'h42 == auto_in_a_bits_source ? count_67 : _GEN_579; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_581 = 9'h43 == auto_in_a_bits_source ? count_68 : _GEN_580; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_582 = 9'h44 == auto_in_a_bits_source ? count_69 : _GEN_581; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_583 = 9'h45 == auto_in_a_bits_source ? count_70 : _GEN_582; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_584 = 9'h46 == auto_in_a_bits_source ? count_71 : _GEN_583; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_585 = 9'h47 == auto_in_a_bits_source ? count_72 : _GEN_584; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_586 = 9'h48 == auto_in_a_bits_source ? count_73 : _GEN_585; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_587 = 9'h49 == auto_in_a_bits_source ? count_74 : _GEN_586; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_588 = 9'h4a == auto_in_a_bits_source ? count_75 : _GEN_587; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_589 = 9'h4b == auto_in_a_bits_source ? count_76 : _GEN_588; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_590 = 9'h4c == auto_in_a_bits_source ? count_77 : _GEN_589; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_591 = 9'h4d == auto_in_a_bits_source ? count_78 : _GEN_590; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_592 = 9'h4e == auto_in_a_bits_source ? count_79 : _GEN_591; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_593 = 9'h4f == auto_in_a_bits_source ? count_80 : _GEN_592; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_594 = 9'h50 == auto_in_a_bits_source ? count_81 : _GEN_593; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_595 = 9'h51 == auto_in_a_bits_source ? count_82 : _GEN_594; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_596 = 9'h52 == auto_in_a_bits_source ? count_83 : _GEN_595; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_597 = 9'h53 == auto_in_a_bits_source ? count_84 : _GEN_596; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_598 = 9'h54 == auto_in_a_bits_source ? count_85 : _GEN_597; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_599 = 9'h55 == auto_in_a_bits_source ? count_86 : _GEN_598; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_600 = 9'h56 == auto_in_a_bits_source ? count_87 : _GEN_599; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_601 = 9'h57 == auto_in_a_bits_source ? count_88 : _GEN_600; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_602 = 9'h58 == auto_in_a_bits_source ? count_89 : _GEN_601; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_603 = 9'h59 == auto_in_a_bits_source ? count_90 : _GEN_602; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_604 = 9'h5a == auto_in_a_bits_source ? count_91 : _GEN_603; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_605 = 9'h5b == auto_in_a_bits_source ? count_92 : _GEN_604; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_606 = 9'h5c == auto_in_a_bits_source ? count_93 : _GEN_605; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_607 = 9'h5d == auto_in_a_bits_source ? count_94 : _GEN_606; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_608 = 9'h5e == auto_in_a_bits_source ? count_95 : _GEN_607; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_609 = 9'h5f == auto_in_a_bits_source ? count_96 : _GEN_608; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_610 = 9'h60 == auto_in_a_bits_source ? count_97 : _GEN_609; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_611 = 9'h61 == auto_in_a_bits_source ? count_98 : _GEN_610; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_612 = 9'h62 == auto_in_a_bits_source ? count_99 : _GEN_611; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_613 = 9'h63 == auto_in_a_bits_source ? count_100 : _GEN_612; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_614 = 9'h64 == auto_in_a_bits_source ? count_101 : _GEN_613; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_615 = 9'h65 == auto_in_a_bits_source ? count_102 : _GEN_614; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_616 = 9'h66 == auto_in_a_bits_source ? count_103 : _GEN_615; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_617 = 9'h67 == auto_in_a_bits_source ? count_104 : _GEN_616; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_618 = 9'h68 == auto_in_a_bits_source ? count_105 : _GEN_617; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_619 = 9'h69 == auto_in_a_bits_source ? count_106 : _GEN_618; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_620 = 9'h6a == auto_in_a_bits_source ? count_107 : _GEN_619; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_621 = 9'h6b == auto_in_a_bits_source ? count_108 : _GEN_620; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_622 = 9'h6c == auto_in_a_bits_source ? count_109 : _GEN_621; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_623 = 9'h6d == auto_in_a_bits_source ? count_110 : _GEN_622; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_624 = 9'h6e == auto_in_a_bits_source ? count_111 : _GEN_623; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_625 = 9'h6f == auto_in_a_bits_source ? count_112 : _GEN_624; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_626 = 9'h70 == auto_in_a_bits_source ? count_113 : _GEN_625; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_627 = 9'h71 == auto_in_a_bits_source ? count_114 : _GEN_626; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_628 = 9'h72 == auto_in_a_bits_source ? count_115 : _GEN_627; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_629 = 9'h73 == auto_in_a_bits_source ? count_116 : _GEN_628; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_630 = 9'h74 == auto_in_a_bits_source ? count_117 : _GEN_629; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_631 = 9'h75 == auto_in_a_bits_source ? count_118 : _GEN_630; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_632 = 9'h76 == auto_in_a_bits_source ? count_119 : _GEN_631; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_633 = 9'h77 == auto_in_a_bits_source ? count_120 : _GEN_632; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_634 = 9'h78 == auto_in_a_bits_source ? count_121 : _GEN_633; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_635 = 9'h79 == auto_in_a_bits_source ? count_122 : _GEN_634; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_636 = 9'h7a == auto_in_a_bits_source ? count_123 : _GEN_635; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_637 = 9'h7b == auto_in_a_bits_source ? count_124 : _GEN_636; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_638 = 9'h7c == auto_in_a_bits_source ? count_125 : _GEN_637; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_639 = 9'h7d == auto_in_a_bits_source ? count_126 : _GEN_638; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_640 = 9'h7e == auto_in_a_bits_source ? count_127 : _GEN_639; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_641 = 9'h7f == auto_in_a_bits_source ? count_128 : _GEN_640; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_642 = 9'h80 == auto_in_a_bits_source ? count_129 : _GEN_641; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_643 = 9'h81 == auto_in_a_bits_source ? count_130 : _GEN_642; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_644 = 9'h82 == auto_in_a_bits_source ? count_131 : _GEN_643; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_645 = 9'h83 == auto_in_a_bits_source ? count_132 : _GEN_644; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_646 = 9'h84 == auto_in_a_bits_source ? count_133 : _GEN_645; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_647 = 9'h85 == auto_in_a_bits_source ? count_134 : _GEN_646; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_648 = 9'h86 == auto_in_a_bits_source ? count_135 : _GEN_647; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_649 = 9'h87 == auto_in_a_bits_source ? count_136 : _GEN_648; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_650 = 9'h88 == auto_in_a_bits_source ? count_137 : _GEN_649; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_651 = 9'h89 == auto_in_a_bits_source ? count_138 : _GEN_650; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_652 = 9'h8a == auto_in_a_bits_source ? count_139 : _GEN_651; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_653 = 9'h8b == auto_in_a_bits_source ? count_140 : _GEN_652; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_654 = 9'h8c == auto_in_a_bits_source ? count_141 : _GEN_653; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_655 = 9'h8d == auto_in_a_bits_source ? count_142 : _GEN_654; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_656 = 9'h8e == auto_in_a_bits_source ? count_143 : _GEN_655; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_657 = 9'h8f == auto_in_a_bits_source ? count_144 : _GEN_656; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_658 = 9'h90 == auto_in_a_bits_source ? count_145 : _GEN_657; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_659 = 9'h91 == auto_in_a_bits_source ? count_146 : _GEN_658; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_660 = 9'h92 == auto_in_a_bits_source ? count_147 : _GEN_659; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_661 = 9'h93 == auto_in_a_bits_source ? count_148 : _GEN_660; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_662 = 9'h94 == auto_in_a_bits_source ? count_149 : _GEN_661; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_663 = 9'h95 == auto_in_a_bits_source ? count_150 : _GEN_662; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_664 = 9'h96 == auto_in_a_bits_source ? count_151 : _GEN_663; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_665 = 9'h97 == auto_in_a_bits_source ? count_152 : _GEN_664; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_666 = 9'h98 == auto_in_a_bits_source ? count_153 : _GEN_665; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_667 = 9'h99 == auto_in_a_bits_source ? count_154 : _GEN_666; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_668 = 9'h9a == auto_in_a_bits_source ? count_155 : _GEN_667; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_669 = 9'h9b == auto_in_a_bits_source ? count_156 : _GEN_668; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_670 = 9'h9c == auto_in_a_bits_source ? count_157 : _GEN_669; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_671 = 9'h9d == auto_in_a_bits_source ? count_158 : _GEN_670; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_672 = 9'h9e == auto_in_a_bits_source ? count_159 : _GEN_671; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_673 = 9'h9f == auto_in_a_bits_source ? count_160 : _GEN_672; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_674 = 9'ha0 == auto_in_a_bits_source ? count_161 : _GEN_673; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_675 = 9'ha1 == auto_in_a_bits_source ? count_162 : _GEN_674; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_676 = 9'ha2 == auto_in_a_bits_source ? count_163 : _GEN_675; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_677 = 9'ha3 == auto_in_a_bits_source ? count_164 : _GEN_676; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_678 = 9'ha4 == auto_in_a_bits_source ? count_165 : _GEN_677; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_679 = 9'ha5 == auto_in_a_bits_source ? count_166 : _GEN_678; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_680 = 9'ha6 == auto_in_a_bits_source ? count_167 : _GEN_679; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_681 = 9'ha7 == auto_in_a_bits_source ? count_168 : _GEN_680; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_682 = 9'ha8 == auto_in_a_bits_source ? count_169 : _GEN_681; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_683 = 9'ha9 == auto_in_a_bits_source ? count_170 : _GEN_682; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_684 = 9'haa == auto_in_a_bits_source ? count_171 : _GEN_683; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_685 = 9'hab == auto_in_a_bits_source ? count_172 : _GEN_684; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_686 = 9'hac == auto_in_a_bits_source ? count_173 : _GEN_685; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_687 = 9'had == auto_in_a_bits_source ? count_174 : _GEN_686; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_688 = 9'hae == auto_in_a_bits_source ? count_175 : _GEN_687; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_689 = 9'haf == auto_in_a_bits_source ? count_176 : _GEN_688; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_690 = 9'hb0 == auto_in_a_bits_source ? count_177 : _GEN_689; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_691 = 9'hb1 == auto_in_a_bits_source ? count_178 : _GEN_690; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_692 = 9'hb2 == auto_in_a_bits_source ? count_179 : _GEN_691; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_693 = 9'hb3 == auto_in_a_bits_source ? count_180 : _GEN_692; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_694 = 9'hb4 == auto_in_a_bits_source ? count_181 : _GEN_693; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_695 = 9'hb5 == auto_in_a_bits_source ? count_182 : _GEN_694; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_696 = 9'hb6 == auto_in_a_bits_source ? count_183 : _GEN_695; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_697 = 9'hb7 == auto_in_a_bits_source ? count_184 : _GEN_696; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_698 = 9'hb8 == auto_in_a_bits_source ? count_185 : _GEN_697; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_699 = 9'hb9 == auto_in_a_bits_source ? count_186 : _GEN_698; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_700 = 9'hba == auto_in_a_bits_source ? count_187 : _GEN_699; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_701 = 9'hbb == auto_in_a_bits_source ? count_188 : _GEN_700; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_702 = 9'hbc == auto_in_a_bits_source ? count_189 : _GEN_701; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_703 = 9'hbd == auto_in_a_bits_source ? count_190 : _GEN_702; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_704 = 9'hbe == auto_in_a_bits_source ? count_191 : _GEN_703; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_705 = 9'hbf == auto_in_a_bits_source ? count_192 : _GEN_704; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_706 = 9'hc0 == auto_in_a_bits_source ? count_193 : _GEN_705; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_707 = 9'hc1 == auto_in_a_bits_source ? count_194 : _GEN_706; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_708 = 9'hc2 == auto_in_a_bits_source ? count_195 : _GEN_707; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_709 = 9'hc3 == auto_in_a_bits_source ? count_196 : _GEN_708; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_710 = 9'hc4 == auto_in_a_bits_source ? count_197 : _GEN_709; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_711 = 9'hc5 == auto_in_a_bits_source ? count_198 : _GEN_710; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_712 = 9'hc6 == auto_in_a_bits_source ? count_199 : _GEN_711; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_713 = 9'hc7 == auto_in_a_bits_source ? count_200 : _GEN_712; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_714 = 9'hc8 == auto_in_a_bits_source ? count_201 : _GEN_713; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_715 = 9'hc9 == auto_in_a_bits_source ? count_202 : _GEN_714; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_716 = 9'hca == auto_in_a_bits_source ? count_203 : _GEN_715; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_717 = 9'hcb == auto_in_a_bits_source ? count_204 : _GEN_716; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_718 = 9'hcc == auto_in_a_bits_source ? count_205 : _GEN_717; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_719 = 9'hcd == auto_in_a_bits_source ? count_206 : _GEN_718; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_720 = 9'hce == auto_in_a_bits_source ? count_207 : _GEN_719; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_721 = 9'hcf == auto_in_a_bits_source ? count_208 : _GEN_720; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_722 = 9'hd0 == auto_in_a_bits_source ? count_209 : _GEN_721; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_723 = 9'hd1 == auto_in_a_bits_source ? count_210 : _GEN_722; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_724 = 9'hd2 == auto_in_a_bits_source ? count_211 : _GEN_723; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_725 = 9'hd3 == auto_in_a_bits_source ? count_212 : _GEN_724; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_726 = 9'hd4 == auto_in_a_bits_source ? count_213 : _GEN_725; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_727 = 9'hd5 == auto_in_a_bits_source ? count_214 : _GEN_726; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_728 = 9'hd6 == auto_in_a_bits_source ? count_215 : _GEN_727; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_729 = 9'hd7 == auto_in_a_bits_source ? count_216 : _GEN_728; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_730 = 9'hd8 == auto_in_a_bits_source ? count_217 : _GEN_729; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_731 = 9'hd9 == auto_in_a_bits_source ? count_218 : _GEN_730; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_732 = 9'hda == auto_in_a_bits_source ? count_219 : _GEN_731; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_733 = 9'hdb == auto_in_a_bits_source ? count_220 : _GEN_732; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_734 = 9'hdc == auto_in_a_bits_source ? count_221 : _GEN_733; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_735 = 9'hdd == auto_in_a_bits_source ? count_222 : _GEN_734; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_736 = 9'hde == auto_in_a_bits_source ? count_223 : _GEN_735; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_737 = 9'hdf == auto_in_a_bits_source ? count_224 : _GEN_736; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_738 = 9'he0 == auto_in_a_bits_source ? count_225 : _GEN_737; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_739 = 9'he1 == auto_in_a_bits_source ? count_226 : _GEN_738; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_740 = 9'he2 == auto_in_a_bits_source ? count_227 : _GEN_739; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_741 = 9'he3 == auto_in_a_bits_source ? count_228 : _GEN_740; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_742 = 9'he4 == auto_in_a_bits_source ? count_229 : _GEN_741; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_743 = 9'he5 == auto_in_a_bits_source ? count_230 : _GEN_742; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_744 = 9'he6 == auto_in_a_bits_source ? count_231 : _GEN_743; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_745 = 9'he7 == auto_in_a_bits_source ? count_232 : _GEN_744; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_746 = 9'he8 == auto_in_a_bits_source ? count_233 : _GEN_745; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_747 = 9'he9 == auto_in_a_bits_source ? count_234 : _GEN_746; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_748 = 9'hea == auto_in_a_bits_source ? count_235 : _GEN_747; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_749 = 9'heb == auto_in_a_bits_source ? count_236 : _GEN_748; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_750 = 9'hec == auto_in_a_bits_source ? count_237 : _GEN_749; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_751 = 9'hed == auto_in_a_bits_source ? count_238 : _GEN_750; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_752 = 9'hee == auto_in_a_bits_source ? count_239 : _GEN_751; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_753 = 9'hef == auto_in_a_bits_source ? count_240 : _GEN_752; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_754 = 9'hf0 == auto_in_a_bits_source ? count_241 : _GEN_753; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_755 = 9'hf1 == auto_in_a_bits_source ? count_242 : _GEN_754; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_756 = 9'hf2 == auto_in_a_bits_source ? count_243 : _GEN_755; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_757 = 9'hf3 == auto_in_a_bits_source ? count_244 : _GEN_756; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_758 = 9'hf4 == auto_in_a_bits_source ? count_245 : _GEN_757; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_759 = 9'hf5 == auto_in_a_bits_source ? count_246 : _GEN_758; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_760 = 9'hf6 == auto_in_a_bits_source ? count_247 : _GEN_759; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_761 = 9'hf7 == auto_in_a_bits_source ? count_248 : _GEN_760; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_762 = 9'hf8 == auto_in_a_bits_source ? count_249 : _GEN_761; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_763 = 9'hf9 == auto_in_a_bits_source ? count_250 : _GEN_762; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_764 = 9'hfa == auto_in_a_bits_source ? count_251 : _GEN_763; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_765 = 9'hfb == auto_in_a_bits_source ? count_252 : _GEN_764; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_766 = 9'hfc == auto_in_a_bits_source ? count_253 : _GEN_765; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_767 = 9'hfd == auto_in_a_bits_source ? count_254 : _GEN_766; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_768 = 9'hfe == auto_in_a_bits_source ? count_255 : _GEN_767; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_769 = 9'hff == auto_in_a_bits_source ? count_256 : _GEN_768; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_770 = 9'h100 == auto_in_a_bits_source ? count_257 : _GEN_769; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_771 = 9'h101 == auto_in_a_bits_source ? count_258 : _GEN_770; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_772 = 9'h102 == auto_in_a_bits_source ? count_259 : _GEN_771; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_773 = 9'h103 == auto_in_a_bits_source ? count_260 : _GEN_772; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_774 = 9'h104 == auto_in_a_bits_source ? count_261 : _GEN_773; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_775 = 9'h105 == auto_in_a_bits_source ? count_262 : _GEN_774; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_776 = 9'h106 == auto_in_a_bits_source ? count_263 : _GEN_775; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_777 = 9'h107 == auto_in_a_bits_source ? count_264 : _GEN_776; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_778 = 9'h108 == auto_in_a_bits_source ? count_265 : _GEN_777; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_779 = 9'h109 == auto_in_a_bits_source ? count_266 : _GEN_778; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_780 = 9'h10a == auto_in_a_bits_source ? count_267 : _GEN_779; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_781 = 9'h10b == auto_in_a_bits_source ? count_268 : _GEN_780; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_782 = 9'h10c == auto_in_a_bits_source ? count_269 : _GEN_781; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_783 = 9'h10d == auto_in_a_bits_source ? count_270 : _GEN_782; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_784 = 9'h10e == auto_in_a_bits_source ? count_271 : _GEN_783; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_785 = 9'h10f == auto_in_a_bits_source ? count_272 : _GEN_784; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_786 = 9'h110 == auto_in_a_bits_source ? count_273 : _GEN_785; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_787 = 9'h111 == auto_in_a_bits_source ? count_274 : _GEN_786; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_788 = 9'h112 == auto_in_a_bits_source ? count_275 : _GEN_787; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_789 = 9'h113 == auto_in_a_bits_source ? count_276 : _GEN_788; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_790 = 9'h114 == auto_in_a_bits_source ? count_277 : _GEN_789; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_791 = 9'h115 == auto_in_a_bits_source ? count_278 : _GEN_790; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_792 = 9'h116 == auto_in_a_bits_source ? count_279 : _GEN_791; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_793 = 9'h117 == auto_in_a_bits_source ? count_280 : _GEN_792; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_794 = 9'h118 == auto_in_a_bits_source ? count_281 : _GEN_793; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_795 = 9'h119 == auto_in_a_bits_source ? count_282 : _GEN_794; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_796 = 9'h11a == auto_in_a_bits_source ? count_283 : _GEN_795; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_797 = 9'h11b == auto_in_a_bits_source ? count_284 : _GEN_796; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_798 = 9'h11c == auto_in_a_bits_source ? count_285 : _GEN_797; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_799 = 9'h11d == auto_in_a_bits_source ? count_286 : _GEN_798; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_800 = 9'h11e == auto_in_a_bits_source ? count_287 : _GEN_799; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_801 = 9'h11f == auto_in_a_bits_source ? count_288 : _GEN_800; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_802 = 9'h120 == auto_in_a_bits_source ? count_289 : _GEN_801; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_803 = 9'h121 == auto_in_a_bits_source ? count_290 : _GEN_802; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_804 = 9'h122 == auto_in_a_bits_source ? count_291 : _GEN_803; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_805 = 9'h123 == auto_in_a_bits_source ? count_292 : _GEN_804; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_806 = 9'h124 == auto_in_a_bits_source ? count_293 : _GEN_805; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_807 = 9'h125 == auto_in_a_bits_source ? count_294 : _GEN_806; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_808 = 9'h126 == auto_in_a_bits_source ? count_295 : _GEN_807; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_809 = 9'h127 == auto_in_a_bits_source ? count_296 : _GEN_808; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_810 = 9'h128 == auto_in_a_bits_source ? count_297 : _GEN_809; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_811 = 9'h129 == auto_in_a_bits_source ? count_298 : _GEN_810; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_812 = 9'h12a == auto_in_a_bits_source ? count_299 : _GEN_811; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_813 = 9'h12b == auto_in_a_bits_source ? count_300 : _GEN_812; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_814 = 9'h12c == auto_in_a_bits_source ? count_301 : _GEN_813; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_815 = 9'h12d == auto_in_a_bits_source ? count_302 : _GEN_814; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_816 = 9'h12e == auto_in_a_bits_source ? count_303 : _GEN_815; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_817 = 9'h12f == auto_in_a_bits_source ? count_304 : _GEN_816; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_818 = 9'h130 == auto_in_a_bits_source ? count_305 : _GEN_817; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_819 = 9'h131 == auto_in_a_bits_source ? count_306 : _GEN_818; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_820 = 9'h132 == auto_in_a_bits_source ? count_307 : _GEN_819; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_821 = 9'h133 == auto_in_a_bits_source ? count_308 : _GEN_820; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_822 = 9'h134 == auto_in_a_bits_source ? count_309 : _GEN_821; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_823 = 9'h135 == auto_in_a_bits_source ? count_310 : _GEN_822; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_824 = 9'h136 == auto_in_a_bits_source ? count_311 : _GEN_823; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_825 = 9'h137 == auto_in_a_bits_source ? count_312 : _GEN_824; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_826 = 9'h138 == auto_in_a_bits_source ? count_313 : _GEN_825; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_827 = 9'h139 == auto_in_a_bits_source ? count_314 : _GEN_826; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_828 = 9'h13a == auto_in_a_bits_source ? count_315 : _GEN_827; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_829 = 9'h13b == auto_in_a_bits_source ? count_316 : _GEN_828; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_830 = 9'h13c == auto_in_a_bits_source ? count_317 : _GEN_829; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_831 = 9'h13d == auto_in_a_bits_source ? count_318 : _GEN_830; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_832 = 9'h13e == auto_in_a_bits_source ? count_319 : _GEN_831; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_833 = 9'h13f == auto_in_a_bits_source ? count_320 : _GEN_832; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_834 = 9'h140 == auto_in_a_bits_source ? count_321 : _GEN_833; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_835 = 9'h141 == auto_in_a_bits_source ? count_322 : _GEN_834; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_836 = 9'h142 == auto_in_a_bits_source ? count_323 : _GEN_835; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_837 = 9'h143 == auto_in_a_bits_source ? count_324 : _GEN_836; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_838 = 9'h144 == auto_in_a_bits_source ? count_325 : _GEN_837; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_839 = 9'h145 == auto_in_a_bits_source ? count_326 : _GEN_838; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_840 = 9'h146 == auto_in_a_bits_source ? count_327 : _GEN_839; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_841 = 9'h147 == auto_in_a_bits_source ? count_328 : _GEN_840; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_842 = 9'h148 == auto_in_a_bits_source ? count_329 : _GEN_841; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_843 = 9'h149 == auto_in_a_bits_source ? count_330 : _GEN_842; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_844 = 9'h14a == auto_in_a_bits_source ? count_331 : _GEN_843; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_845 = 9'h14b == auto_in_a_bits_source ? count_332 : _GEN_844; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_846 = 9'h14c == auto_in_a_bits_source ? count_333 : _GEN_845; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_847 = 9'h14d == auto_in_a_bits_source ? count_334 : _GEN_846; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_848 = 9'h14e == auto_in_a_bits_source ? count_335 : _GEN_847; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_849 = 9'h14f == auto_in_a_bits_source ? count_336 : _GEN_848; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_850 = 9'h150 == auto_in_a_bits_source ? count_337 : _GEN_849; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_851 = 9'h151 == auto_in_a_bits_source ? count_338 : _GEN_850; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_852 = 9'h152 == auto_in_a_bits_source ? count_339 : _GEN_851; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_853 = 9'h153 == auto_in_a_bits_source ? count_340 : _GEN_852; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_854 = 9'h154 == auto_in_a_bits_source ? count_341 : _GEN_853; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_855 = 9'h155 == auto_in_a_bits_source ? count_342 : _GEN_854; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_856 = 9'h156 == auto_in_a_bits_source ? count_343 : _GEN_855; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_857 = 9'h157 == auto_in_a_bits_source ? count_344 : _GEN_856; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_858 = 9'h158 == auto_in_a_bits_source ? count_345 : _GEN_857; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_859 = 9'h159 == auto_in_a_bits_source ? count_346 : _GEN_858; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_860 = 9'h15a == auto_in_a_bits_source ? count_347 : _GEN_859; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_861 = 9'h15b == auto_in_a_bits_source ? count_348 : _GEN_860; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_862 = 9'h15c == auto_in_a_bits_source ? count_349 : _GEN_861; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_863 = 9'h15d == auto_in_a_bits_source ? count_350 : _GEN_862; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_864 = 9'h15e == auto_in_a_bits_source ? count_351 : _GEN_863; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_865 = 9'h15f == auto_in_a_bits_source ? count_352 : _GEN_864; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_866 = 9'h160 == auto_in_a_bits_source ? count_353 : _GEN_865; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_867 = 9'h161 == auto_in_a_bits_source ? count_354 : _GEN_866; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_868 = 9'h162 == auto_in_a_bits_source ? count_355 : _GEN_867; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_869 = 9'h163 == auto_in_a_bits_source ? count_356 : _GEN_868; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_870 = 9'h164 == auto_in_a_bits_source ? count_357 : _GEN_869; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_871 = 9'h165 == auto_in_a_bits_source ? count_358 : _GEN_870; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_872 = 9'h166 == auto_in_a_bits_source ? count_359 : _GEN_871; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_873 = 9'h167 == auto_in_a_bits_source ? count_360 : _GEN_872; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_874 = 9'h168 == auto_in_a_bits_source ? count_361 : _GEN_873; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_875 = 9'h169 == auto_in_a_bits_source ? count_362 : _GEN_874; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_876 = 9'h16a == auto_in_a_bits_source ? count_363 : _GEN_875; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_877 = 9'h16b == auto_in_a_bits_source ? count_364 : _GEN_876; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_878 = 9'h16c == auto_in_a_bits_source ? count_365 : _GEN_877; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_879 = 9'h16d == auto_in_a_bits_source ? count_366 : _GEN_878; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_880 = 9'h16e == auto_in_a_bits_source ? count_367 : _GEN_879; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_881 = 9'h16f == auto_in_a_bits_source ? count_368 : _GEN_880; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_882 = 9'h170 == auto_in_a_bits_source ? count_369 : _GEN_881; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_883 = 9'h171 == auto_in_a_bits_source ? count_370 : _GEN_882; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_884 = 9'h172 == auto_in_a_bits_source ? count_371 : _GEN_883; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_885 = 9'h173 == auto_in_a_bits_source ? count_372 : _GEN_884; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_886 = 9'h174 == auto_in_a_bits_source ? count_373 : _GEN_885; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_887 = 9'h175 == auto_in_a_bits_source ? count_374 : _GEN_886; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_888 = 9'h176 == auto_in_a_bits_source ? count_375 : _GEN_887; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_889 = 9'h177 == auto_in_a_bits_source ? count_376 : _GEN_888; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_890 = 9'h178 == auto_in_a_bits_source ? count_377 : _GEN_889; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_891 = 9'h179 == auto_in_a_bits_source ? count_378 : _GEN_890; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_892 = 9'h17a == auto_in_a_bits_source ? count_379 : _GEN_891; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_893 = 9'h17b == auto_in_a_bits_source ? count_380 : _GEN_892; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_894 = 9'h17c == auto_in_a_bits_source ? count_381 : _GEN_893; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_895 = 9'h17d == auto_in_a_bits_source ? count_382 : _GEN_894; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_896 = 9'h17e == auto_in_a_bits_source ? count_383 : _GEN_895; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_897 = 9'h17f == auto_in_a_bits_source ? count_384 : _GEN_896; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_898 = 9'h180 == auto_in_a_bits_source ? count_385 : _GEN_897; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_899 = 9'h181 == auto_in_a_bits_source ? count_386 : _GEN_898; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_900 = 9'h182 == auto_in_a_bits_source ? count_387 : _GEN_899; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_901 = 9'h183 == auto_in_a_bits_source ? count_388 : _GEN_900; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_902 = 9'h184 == auto_in_a_bits_source ? count_389 : _GEN_901; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_903 = 9'h185 == auto_in_a_bits_source ? count_390 : _GEN_902; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_904 = 9'h186 == auto_in_a_bits_source ? count_391 : _GEN_903; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_905 = 9'h187 == auto_in_a_bits_source ? count_392 : _GEN_904; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_906 = 9'h188 == auto_in_a_bits_source ? count_393 : _GEN_905; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_907 = 9'h189 == auto_in_a_bits_source ? count_394 : _GEN_906; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_908 = 9'h18a == auto_in_a_bits_source ? count_395 : _GEN_907; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_909 = 9'h18b == auto_in_a_bits_source ? count_396 : _GEN_908; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_910 = 9'h18c == auto_in_a_bits_source ? count_397 : _GEN_909; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_911 = 9'h18d == auto_in_a_bits_source ? count_398 : _GEN_910; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_912 = 9'h18e == auto_in_a_bits_source ? count_399 : _GEN_911; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_913 = 9'h18f == auto_in_a_bits_source ? count_400 : _GEN_912; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_914 = 9'h190 == auto_in_a_bits_source ? count_401 : _GEN_913; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_915 = 9'h191 == auto_in_a_bits_source ? count_402 : _GEN_914; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_916 = 9'h192 == auto_in_a_bits_source ? count_403 : _GEN_915; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_917 = 9'h193 == auto_in_a_bits_source ? count_404 : _GEN_916; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_918 = 9'h194 == auto_in_a_bits_source ? count_405 : _GEN_917; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_919 = 9'h195 == auto_in_a_bits_source ? count_406 : _GEN_918; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_920 = 9'h196 == auto_in_a_bits_source ? count_407 : _GEN_919; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_921 = 9'h197 == auto_in_a_bits_source ? count_408 : _GEN_920; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_922 = 9'h198 == auto_in_a_bits_source ? count_409 : _GEN_921; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_923 = 9'h199 == auto_in_a_bits_source ? count_410 : _GEN_922; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_924 = 9'h19a == auto_in_a_bits_source ? count_411 : _GEN_923; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_925 = 9'h19b == auto_in_a_bits_source ? count_412 : _GEN_924; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_926 = 9'h19c == auto_in_a_bits_source ? count_413 : _GEN_925; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_927 = 9'h19d == auto_in_a_bits_source ? count_414 : _GEN_926; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_928 = 9'h19e == auto_in_a_bits_source ? count_415 : _GEN_927; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_929 = 9'h19f == auto_in_a_bits_source ? count_416 : _GEN_928; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_930 = 9'h1a0 == auto_in_a_bits_source ? count_417 : _GEN_929; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_931 = 9'h1a1 == auto_in_a_bits_source ? count_418 : _GEN_930; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_932 = 9'h1a2 == auto_in_a_bits_source ? count_419 : _GEN_931; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_933 = 9'h1a3 == auto_in_a_bits_source ? count_420 : _GEN_932; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_934 = 9'h1a4 == auto_in_a_bits_source ? count_421 : _GEN_933; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_935 = 9'h1a5 == auto_in_a_bits_source ? count_422 : _GEN_934; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_936 = 9'h1a6 == auto_in_a_bits_source ? count_423 : _GEN_935; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_937 = 9'h1a7 == auto_in_a_bits_source ? count_424 : _GEN_936; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_938 = 9'h1a8 == auto_in_a_bits_source ? count_425 : _GEN_937; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_939 = 9'h1a9 == auto_in_a_bits_source ? count_426 : _GEN_938; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_940 = 9'h1aa == auto_in_a_bits_source ? count_427 : _GEN_939; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_941 = 9'h1ab == auto_in_a_bits_source ? count_428 : _GEN_940; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_942 = 9'h1ac == auto_in_a_bits_source ? count_429 : _GEN_941; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_943 = 9'h1ad == auto_in_a_bits_source ? count_430 : _GEN_942; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_944 = 9'h1ae == auto_in_a_bits_source ? count_431 : _GEN_943; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_945 = 9'h1af == auto_in_a_bits_source ? count_432 : _GEN_944; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_946 = 9'h1b0 == auto_in_a_bits_source ? count_433 : _GEN_945; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_947 = 9'h1b1 == auto_in_a_bits_source ? count_434 : _GEN_946; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_948 = 9'h1b2 == auto_in_a_bits_source ? count_435 : _GEN_947; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_949 = 9'h1b3 == auto_in_a_bits_source ? count_436 : _GEN_948; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_950 = 9'h1b4 == auto_in_a_bits_source ? count_437 : _GEN_949; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_951 = 9'h1b5 == auto_in_a_bits_source ? count_438 : _GEN_950; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_952 = 9'h1b6 == auto_in_a_bits_source ? count_439 : _GEN_951; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_953 = 9'h1b7 == auto_in_a_bits_source ? count_440 : _GEN_952; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_954 = 9'h1b8 == auto_in_a_bits_source ? count_441 : _GEN_953; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_955 = 9'h1b9 == auto_in_a_bits_source ? count_442 : _GEN_954; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_956 = 9'h1ba == auto_in_a_bits_source ? count_443 : _GEN_955; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_957 = 9'h1bb == auto_in_a_bits_source ? count_444 : _GEN_956; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_958 = 9'h1bc == auto_in_a_bits_source ? count_445 : _GEN_957; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_959 = 9'h1bd == auto_in_a_bits_source ? count_446 : _GEN_958; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_960 = 9'h1be == auto_in_a_bits_source ? count_447 : _GEN_959; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_961 = 9'h1bf == auto_in_a_bits_source ? count_448 : _GEN_960; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_962 = 9'h1c0 == auto_in_a_bits_source ? count_449 : _GEN_961; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_963 = 9'h1c1 == auto_in_a_bits_source ? count_450 : _GEN_962; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_964 = 9'h1c2 == auto_in_a_bits_source ? count_451 : _GEN_963; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_965 = 9'h1c3 == auto_in_a_bits_source ? count_452 : _GEN_964; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_966 = 9'h1c4 == auto_in_a_bits_source ? count_453 : _GEN_965; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_967 = 9'h1c5 == auto_in_a_bits_source ? count_454 : _GEN_966; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_968 = 9'h1c6 == auto_in_a_bits_source ? count_455 : _GEN_967; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_969 = 9'h1c7 == auto_in_a_bits_source ? count_456 : _GEN_968; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_970 = 9'h1c8 == auto_in_a_bits_source ? count_457 : _GEN_969; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_971 = 9'h1c9 == auto_in_a_bits_source ? count_458 : _GEN_970; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_972 = 9'h1ca == auto_in_a_bits_source ? count_459 : _GEN_971; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_973 = 9'h1cb == auto_in_a_bits_source ? count_460 : _GEN_972; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_974 = 9'h1cc == auto_in_a_bits_source ? count_461 : _GEN_973; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_975 = 9'h1cd == auto_in_a_bits_source ? count_462 : _GEN_974; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_976 = 9'h1ce == auto_in_a_bits_source ? count_463 : _GEN_975; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_977 = 9'h1cf == auto_in_a_bits_source ? count_464 : _GEN_976; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_978 = 9'h1d0 == auto_in_a_bits_source ? count_465 : _GEN_977; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_979 = 9'h1d1 == auto_in_a_bits_source ? count_466 : _GEN_978; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_980 = 9'h1d2 == auto_in_a_bits_source ? count_467 : _GEN_979; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_981 = 9'h1d3 == auto_in_a_bits_source ? count_468 : _GEN_980; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_982 = 9'h1d4 == auto_in_a_bits_source ? count_469 : _GEN_981; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_983 = 9'h1d5 == auto_in_a_bits_source ? count_470 : _GEN_982; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_984 = 9'h1d6 == auto_in_a_bits_source ? count_471 : _GEN_983; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_985 = 9'h1d7 == auto_in_a_bits_source ? count_472 : _GEN_984; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_986 = 9'h1d8 == auto_in_a_bits_source ? count_473 : _GEN_985; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_987 = 9'h1d9 == auto_in_a_bits_source ? count_474 : _GEN_986; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_988 = 9'h1da == auto_in_a_bits_source ? count_475 : _GEN_987; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_989 = 9'h1db == auto_in_a_bits_source ? count_476 : _GEN_988; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_990 = 9'h1dc == auto_in_a_bits_source ? count_477 : _GEN_989; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_991 = 9'h1dd == auto_in_a_bits_source ? count_478 : _GEN_990; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_992 = 9'h1de == auto_in_a_bits_source ? count_479 : _GEN_991; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_993 = 9'h1df == auto_in_a_bits_source ? count_480 : _GEN_992; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_994 = 9'h1e0 == auto_in_a_bits_source ? count_481 : _GEN_993; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_995 = 9'h1e1 == auto_in_a_bits_source ? count_482 : _GEN_994; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_996 = 9'h1e2 == auto_in_a_bits_source ? count_483 : _GEN_995; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_997 = 9'h1e3 == auto_in_a_bits_source ? count_484 : _GEN_996; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_998 = 9'h1e4 == auto_in_a_bits_source ? count_485 : _GEN_997; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_999 = 9'h1e5 == auto_in_a_bits_source ? count_486 : _GEN_998; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1000 = 9'h1e6 == auto_in_a_bits_source ? count_487 : _GEN_999; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1001 = 9'h1e7 == auto_in_a_bits_source ? count_488 : _GEN_1000; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1002 = 9'h1e8 == auto_in_a_bits_source ? count_489 : _GEN_1001; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1003 = 9'h1e9 == auto_in_a_bits_source ? count_490 : _GEN_1002; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1004 = 9'h1ea == auto_in_a_bits_source ? count_491 : _GEN_1003; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1005 = 9'h1eb == auto_in_a_bits_source ? count_492 : _GEN_1004; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1006 = 9'h1ec == auto_in_a_bits_source ? count_493 : _GEN_1005; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1007 = 9'h1ed == auto_in_a_bits_source ? count_494 : _GEN_1006; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1008 = 9'h1ee == auto_in_a_bits_source ? count_495 : _GEN_1007; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1009 = 9'h1ef == auto_in_a_bits_source ? count_496 : _GEN_1008; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1010 = 9'h1f0 == auto_in_a_bits_source ? count_497 : _GEN_1009; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1011 = 9'h1f1 == auto_in_a_bits_source ? count_498 : _GEN_1010; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1012 = 9'h1f2 == auto_in_a_bits_source ? count_499 : _GEN_1011; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1013 = 9'h1f3 == auto_in_a_bits_source ? count_500 : _GEN_1012; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1014 = 9'h1f4 == auto_in_a_bits_source ? count_501 : _GEN_1013; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1015 = 9'h1f5 == auto_in_a_bits_source ? count_502 : _GEN_1014; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1016 = 9'h1f6 == auto_in_a_bits_source ? count_503 : _GEN_1015; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1017 = 9'h1f7 == auto_in_a_bits_source ? count_504 : _GEN_1016; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1018 = 9'h1f8 == auto_in_a_bits_source ? count_505 : _GEN_1017; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1019 = 9'h1f9 == auto_in_a_bits_source ? count_506 : _GEN_1018; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1020 = 9'h1fa == auto_in_a_bits_source ? count_507 : _GEN_1019; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1021 = 9'h1fb == auto_in_a_bits_source ? count_508 : _GEN_1020; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1022 = 9'h1fc == auto_in_a_bits_source ? count_509 : _GEN_1021; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1023 = 9'h1fd == auto_in_a_bits_source ? count_510 : _GEN_1022; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1024 = 9'h1fe == auto_in_a_bits_source ? count_511 : _GEN_1023; // @[ToAXI4.scala 195:{49,49}]
  wire  _GEN_1025 = 9'h1ff == auto_in_a_bits_source ? count_512 : _GEN_1024; // @[ToAXI4.scala 195:{49,49}]
  reg [2:0] counter; // @[Edges.scala 228:27]
  wire  a_first = counter == 3'h0; // @[Edges.scala 230:25]
  wire  stall = _GEN_1025 & a_first; // @[ToAXI4.scala 195:49]
  wire  _bundleIn_0_a_ready_T = ~stall; // @[ToAXI4.scala 196:21]
  reg  doneAW; // @[ToAXI4.scala 161:30]
  wire  out_arw_ready = queue_arw_deq_io_enq_ready; // @[ToAXI4.scala 147:25 Decoupled.scala 365:17]
  wire  _bundleIn_0_a_ready_T_1 = doneAW | out_arw_ready; // @[ToAXI4.scala 196:52]
  wire  out_w_ready = deq_io_enq_ready; // @[ToAXI4.scala 148:23 Decoupled.scala 365:17]
  wire  _bundleIn_0_a_ready_T_3 = a_isPut ? (doneAW | out_arw_ready) & out_w_ready : out_arw_ready; // @[ToAXI4.scala 196:34]
  wire  bundleIn_0_a_ready = ~stall & _bundleIn_0_a_ready_T_3; // @[ToAXI4.scala 196:28]
  wire  _T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 50:35]
  wire [12:0] _beats1_decode_T_1 = 13'h3f << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] beats1_decode = _beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire [2:0] beats1 = a_isPut ? beats1_decode : 3'h0; // @[Edges.scala 220:14]
  wire [2:0] counter1 = counter - 3'h1; // @[Edges.scala 229:28]
  wire  a_last = counter == 3'h1 | beats1 == 3'h0; // @[Edges.scala 231:37]
  wire  queue_arw_bits_wen = queue_arw_deq_io_deq_bits_wen; // @[Decoupled.scala 401:19 402:14]
  wire  queue_arw_valid = queue_arw_deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  wire [8:0] _GEN_3 = 9'h1 == auto_in_a_bits_source ? 9'h1 : 9'h0; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_4 = 9'h2 == auto_in_a_bits_source ? 9'h2 : _GEN_3; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_5 = 9'h3 == auto_in_a_bits_source ? 9'h3 : _GEN_4; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_6 = 9'h4 == auto_in_a_bits_source ? 9'h4 : _GEN_5; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_7 = 9'h5 == auto_in_a_bits_source ? 9'h5 : _GEN_6; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_8 = 9'h6 == auto_in_a_bits_source ? 9'h6 : _GEN_7; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_9 = 9'h7 == auto_in_a_bits_source ? 9'h7 : _GEN_8; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_10 = 9'h8 == auto_in_a_bits_source ? 9'h8 : _GEN_9; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_11 = 9'h9 == auto_in_a_bits_source ? 9'h9 : _GEN_10; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_12 = 9'ha == auto_in_a_bits_source ? 9'ha : _GEN_11; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_13 = 9'hb == auto_in_a_bits_source ? 9'hb : _GEN_12; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_14 = 9'hc == auto_in_a_bits_source ? 9'hc : _GEN_13; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_15 = 9'hd == auto_in_a_bits_source ? 9'hd : _GEN_14; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_16 = 9'he == auto_in_a_bits_source ? 9'he : _GEN_15; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_17 = 9'hf == auto_in_a_bits_source ? 9'hf : _GEN_16; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_18 = 9'h10 == auto_in_a_bits_source ? 9'h10 : _GEN_17; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_19 = 9'h11 == auto_in_a_bits_source ? 9'h11 : _GEN_18; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_20 = 9'h12 == auto_in_a_bits_source ? 9'h12 : _GEN_19; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_21 = 9'h13 == auto_in_a_bits_source ? 9'h13 : _GEN_20; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_22 = 9'h14 == auto_in_a_bits_source ? 9'h14 : _GEN_21; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_23 = 9'h15 == auto_in_a_bits_source ? 9'h15 : _GEN_22; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_24 = 9'h16 == auto_in_a_bits_source ? 9'h16 : _GEN_23; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_25 = 9'h17 == auto_in_a_bits_source ? 9'h17 : _GEN_24; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_26 = 9'h18 == auto_in_a_bits_source ? 9'h18 : _GEN_25; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_27 = 9'h19 == auto_in_a_bits_source ? 9'h19 : _GEN_26; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_28 = 9'h1a == auto_in_a_bits_source ? 9'h1a : _GEN_27; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_29 = 9'h1b == auto_in_a_bits_source ? 9'h1b : _GEN_28; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_30 = 9'h1c == auto_in_a_bits_source ? 9'h1c : _GEN_29; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_31 = 9'h1d == auto_in_a_bits_source ? 9'h1d : _GEN_30; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_32 = 9'h1e == auto_in_a_bits_source ? 9'h1e : _GEN_31; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_33 = 9'h1f == auto_in_a_bits_source ? 9'h1f : _GEN_32; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_34 = 9'h20 == auto_in_a_bits_source ? 9'h20 : _GEN_33; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_35 = 9'h21 == auto_in_a_bits_source ? 9'h21 : _GEN_34; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_36 = 9'h22 == auto_in_a_bits_source ? 9'h22 : _GEN_35; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_37 = 9'h23 == auto_in_a_bits_source ? 9'h23 : _GEN_36; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_38 = 9'h24 == auto_in_a_bits_source ? 9'h24 : _GEN_37; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_39 = 9'h25 == auto_in_a_bits_source ? 9'h25 : _GEN_38; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_40 = 9'h26 == auto_in_a_bits_source ? 9'h26 : _GEN_39; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_41 = 9'h27 == auto_in_a_bits_source ? 9'h27 : _GEN_40; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_42 = 9'h28 == auto_in_a_bits_source ? 9'h28 : _GEN_41; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_43 = 9'h29 == auto_in_a_bits_source ? 9'h29 : _GEN_42; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_44 = 9'h2a == auto_in_a_bits_source ? 9'h2a : _GEN_43; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_45 = 9'h2b == auto_in_a_bits_source ? 9'h2b : _GEN_44; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_46 = 9'h2c == auto_in_a_bits_source ? 9'h2c : _GEN_45; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_47 = 9'h2d == auto_in_a_bits_source ? 9'h2d : _GEN_46; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_48 = 9'h2e == auto_in_a_bits_source ? 9'h2e : _GEN_47; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_49 = 9'h2f == auto_in_a_bits_source ? 9'h2f : _GEN_48; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_50 = 9'h30 == auto_in_a_bits_source ? 9'h30 : _GEN_49; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_51 = 9'h31 == auto_in_a_bits_source ? 9'h31 : _GEN_50; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_52 = 9'h32 == auto_in_a_bits_source ? 9'h32 : _GEN_51; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_53 = 9'h33 == auto_in_a_bits_source ? 9'h33 : _GEN_52; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_54 = 9'h34 == auto_in_a_bits_source ? 9'h34 : _GEN_53; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_55 = 9'h35 == auto_in_a_bits_source ? 9'h35 : _GEN_54; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_56 = 9'h36 == auto_in_a_bits_source ? 9'h36 : _GEN_55; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_57 = 9'h37 == auto_in_a_bits_source ? 9'h37 : _GEN_56; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_58 = 9'h38 == auto_in_a_bits_source ? 9'h38 : _GEN_57; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_59 = 9'h39 == auto_in_a_bits_source ? 9'h39 : _GEN_58; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_60 = 9'h3a == auto_in_a_bits_source ? 9'h3a : _GEN_59; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_61 = 9'h3b == auto_in_a_bits_source ? 9'h3b : _GEN_60; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_62 = 9'h3c == auto_in_a_bits_source ? 9'h3c : _GEN_61; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_63 = 9'h3d == auto_in_a_bits_source ? 9'h3d : _GEN_62; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_64 = 9'h3e == auto_in_a_bits_source ? 9'h3e : _GEN_63; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_65 = 9'h3f == auto_in_a_bits_source ? 9'h3f : _GEN_64; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_66 = 9'h40 == auto_in_a_bits_source ? 9'h40 : _GEN_65; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_67 = 9'h41 == auto_in_a_bits_source ? 9'h41 : _GEN_66; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_68 = 9'h42 == auto_in_a_bits_source ? 9'h42 : _GEN_67; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_69 = 9'h43 == auto_in_a_bits_source ? 9'h43 : _GEN_68; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_70 = 9'h44 == auto_in_a_bits_source ? 9'h44 : _GEN_69; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_71 = 9'h45 == auto_in_a_bits_source ? 9'h45 : _GEN_70; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_72 = 9'h46 == auto_in_a_bits_source ? 9'h46 : _GEN_71; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_73 = 9'h47 == auto_in_a_bits_source ? 9'h47 : _GEN_72; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_74 = 9'h48 == auto_in_a_bits_source ? 9'h48 : _GEN_73; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_75 = 9'h49 == auto_in_a_bits_source ? 9'h49 : _GEN_74; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_76 = 9'h4a == auto_in_a_bits_source ? 9'h4a : _GEN_75; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_77 = 9'h4b == auto_in_a_bits_source ? 9'h4b : _GEN_76; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_78 = 9'h4c == auto_in_a_bits_source ? 9'h4c : _GEN_77; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_79 = 9'h4d == auto_in_a_bits_source ? 9'h4d : _GEN_78; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_80 = 9'h4e == auto_in_a_bits_source ? 9'h4e : _GEN_79; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_81 = 9'h4f == auto_in_a_bits_source ? 9'h4f : _GEN_80; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_82 = 9'h50 == auto_in_a_bits_source ? 9'h50 : _GEN_81; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_83 = 9'h51 == auto_in_a_bits_source ? 9'h51 : _GEN_82; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_84 = 9'h52 == auto_in_a_bits_source ? 9'h52 : _GEN_83; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_85 = 9'h53 == auto_in_a_bits_source ? 9'h53 : _GEN_84; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_86 = 9'h54 == auto_in_a_bits_source ? 9'h54 : _GEN_85; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_87 = 9'h55 == auto_in_a_bits_source ? 9'h55 : _GEN_86; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_88 = 9'h56 == auto_in_a_bits_source ? 9'h56 : _GEN_87; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_89 = 9'h57 == auto_in_a_bits_source ? 9'h57 : _GEN_88; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_90 = 9'h58 == auto_in_a_bits_source ? 9'h58 : _GEN_89; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_91 = 9'h59 == auto_in_a_bits_source ? 9'h59 : _GEN_90; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_92 = 9'h5a == auto_in_a_bits_source ? 9'h5a : _GEN_91; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_93 = 9'h5b == auto_in_a_bits_source ? 9'h5b : _GEN_92; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_94 = 9'h5c == auto_in_a_bits_source ? 9'h5c : _GEN_93; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_95 = 9'h5d == auto_in_a_bits_source ? 9'h5d : _GEN_94; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_96 = 9'h5e == auto_in_a_bits_source ? 9'h5e : _GEN_95; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_97 = 9'h5f == auto_in_a_bits_source ? 9'h5f : _GEN_96; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_98 = 9'h60 == auto_in_a_bits_source ? 9'h60 : _GEN_97; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_99 = 9'h61 == auto_in_a_bits_source ? 9'h61 : _GEN_98; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_100 = 9'h62 == auto_in_a_bits_source ? 9'h62 : _GEN_99; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_101 = 9'h63 == auto_in_a_bits_source ? 9'h63 : _GEN_100; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_102 = 9'h64 == auto_in_a_bits_source ? 9'h64 : _GEN_101; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_103 = 9'h65 == auto_in_a_bits_source ? 9'h65 : _GEN_102; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_104 = 9'h66 == auto_in_a_bits_source ? 9'h66 : _GEN_103; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_105 = 9'h67 == auto_in_a_bits_source ? 9'h67 : _GEN_104; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_106 = 9'h68 == auto_in_a_bits_source ? 9'h68 : _GEN_105; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_107 = 9'h69 == auto_in_a_bits_source ? 9'h69 : _GEN_106; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_108 = 9'h6a == auto_in_a_bits_source ? 9'h6a : _GEN_107; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_109 = 9'h6b == auto_in_a_bits_source ? 9'h6b : _GEN_108; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_110 = 9'h6c == auto_in_a_bits_source ? 9'h6c : _GEN_109; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_111 = 9'h6d == auto_in_a_bits_source ? 9'h6d : _GEN_110; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_112 = 9'h6e == auto_in_a_bits_source ? 9'h6e : _GEN_111; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_113 = 9'h6f == auto_in_a_bits_source ? 9'h6f : _GEN_112; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_114 = 9'h70 == auto_in_a_bits_source ? 9'h70 : _GEN_113; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_115 = 9'h71 == auto_in_a_bits_source ? 9'h71 : _GEN_114; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_116 = 9'h72 == auto_in_a_bits_source ? 9'h72 : _GEN_115; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_117 = 9'h73 == auto_in_a_bits_source ? 9'h73 : _GEN_116; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_118 = 9'h74 == auto_in_a_bits_source ? 9'h74 : _GEN_117; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_119 = 9'h75 == auto_in_a_bits_source ? 9'h75 : _GEN_118; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_120 = 9'h76 == auto_in_a_bits_source ? 9'h76 : _GEN_119; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_121 = 9'h77 == auto_in_a_bits_source ? 9'h77 : _GEN_120; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_122 = 9'h78 == auto_in_a_bits_source ? 9'h78 : _GEN_121; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_123 = 9'h79 == auto_in_a_bits_source ? 9'h79 : _GEN_122; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_124 = 9'h7a == auto_in_a_bits_source ? 9'h7a : _GEN_123; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_125 = 9'h7b == auto_in_a_bits_source ? 9'h7b : _GEN_124; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_126 = 9'h7c == auto_in_a_bits_source ? 9'h7c : _GEN_125; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_127 = 9'h7d == auto_in_a_bits_source ? 9'h7d : _GEN_126; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_128 = 9'h7e == auto_in_a_bits_source ? 9'h7e : _GEN_127; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_129 = 9'h7f == auto_in_a_bits_source ? 9'h7f : _GEN_128; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_130 = 9'h80 == auto_in_a_bits_source ? 9'h80 : _GEN_129; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_131 = 9'h81 == auto_in_a_bits_source ? 9'h81 : _GEN_130; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_132 = 9'h82 == auto_in_a_bits_source ? 9'h82 : _GEN_131; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_133 = 9'h83 == auto_in_a_bits_source ? 9'h83 : _GEN_132; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_134 = 9'h84 == auto_in_a_bits_source ? 9'h84 : _GEN_133; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_135 = 9'h85 == auto_in_a_bits_source ? 9'h85 : _GEN_134; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_136 = 9'h86 == auto_in_a_bits_source ? 9'h86 : _GEN_135; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_137 = 9'h87 == auto_in_a_bits_source ? 9'h87 : _GEN_136; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_138 = 9'h88 == auto_in_a_bits_source ? 9'h88 : _GEN_137; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_139 = 9'h89 == auto_in_a_bits_source ? 9'h89 : _GEN_138; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_140 = 9'h8a == auto_in_a_bits_source ? 9'h8a : _GEN_139; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_141 = 9'h8b == auto_in_a_bits_source ? 9'h8b : _GEN_140; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_142 = 9'h8c == auto_in_a_bits_source ? 9'h8c : _GEN_141; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_143 = 9'h8d == auto_in_a_bits_source ? 9'h8d : _GEN_142; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_144 = 9'h8e == auto_in_a_bits_source ? 9'h8e : _GEN_143; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_145 = 9'h8f == auto_in_a_bits_source ? 9'h8f : _GEN_144; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_146 = 9'h90 == auto_in_a_bits_source ? 9'h90 : _GEN_145; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_147 = 9'h91 == auto_in_a_bits_source ? 9'h91 : _GEN_146; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_148 = 9'h92 == auto_in_a_bits_source ? 9'h92 : _GEN_147; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_149 = 9'h93 == auto_in_a_bits_source ? 9'h93 : _GEN_148; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_150 = 9'h94 == auto_in_a_bits_source ? 9'h94 : _GEN_149; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_151 = 9'h95 == auto_in_a_bits_source ? 9'h95 : _GEN_150; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_152 = 9'h96 == auto_in_a_bits_source ? 9'h96 : _GEN_151; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_153 = 9'h97 == auto_in_a_bits_source ? 9'h97 : _GEN_152; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_154 = 9'h98 == auto_in_a_bits_source ? 9'h98 : _GEN_153; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_155 = 9'h99 == auto_in_a_bits_source ? 9'h99 : _GEN_154; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_156 = 9'h9a == auto_in_a_bits_source ? 9'h9a : _GEN_155; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_157 = 9'h9b == auto_in_a_bits_source ? 9'h9b : _GEN_156; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_158 = 9'h9c == auto_in_a_bits_source ? 9'h9c : _GEN_157; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_159 = 9'h9d == auto_in_a_bits_source ? 9'h9d : _GEN_158; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_160 = 9'h9e == auto_in_a_bits_source ? 9'h9e : _GEN_159; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_161 = 9'h9f == auto_in_a_bits_source ? 9'h9f : _GEN_160; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_162 = 9'ha0 == auto_in_a_bits_source ? 9'ha0 : _GEN_161; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_163 = 9'ha1 == auto_in_a_bits_source ? 9'ha1 : _GEN_162; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_164 = 9'ha2 == auto_in_a_bits_source ? 9'ha2 : _GEN_163; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_165 = 9'ha3 == auto_in_a_bits_source ? 9'ha3 : _GEN_164; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_166 = 9'ha4 == auto_in_a_bits_source ? 9'ha4 : _GEN_165; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_167 = 9'ha5 == auto_in_a_bits_source ? 9'ha5 : _GEN_166; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_168 = 9'ha6 == auto_in_a_bits_source ? 9'ha6 : _GEN_167; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_169 = 9'ha7 == auto_in_a_bits_source ? 9'ha7 : _GEN_168; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_170 = 9'ha8 == auto_in_a_bits_source ? 9'ha8 : _GEN_169; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_171 = 9'ha9 == auto_in_a_bits_source ? 9'ha9 : _GEN_170; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_172 = 9'haa == auto_in_a_bits_source ? 9'haa : _GEN_171; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_173 = 9'hab == auto_in_a_bits_source ? 9'hab : _GEN_172; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_174 = 9'hac == auto_in_a_bits_source ? 9'hac : _GEN_173; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_175 = 9'had == auto_in_a_bits_source ? 9'had : _GEN_174; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_176 = 9'hae == auto_in_a_bits_source ? 9'hae : _GEN_175; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_177 = 9'haf == auto_in_a_bits_source ? 9'haf : _GEN_176; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_178 = 9'hb0 == auto_in_a_bits_source ? 9'hb0 : _GEN_177; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_179 = 9'hb1 == auto_in_a_bits_source ? 9'hb1 : _GEN_178; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_180 = 9'hb2 == auto_in_a_bits_source ? 9'hb2 : _GEN_179; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_181 = 9'hb3 == auto_in_a_bits_source ? 9'hb3 : _GEN_180; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_182 = 9'hb4 == auto_in_a_bits_source ? 9'hb4 : _GEN_181; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_183 = 9'hb5 == auto_in_a_bits_source ? 9'hb5 : _GEN_182; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_184 = 9'hb6 == auto_in_a_bits_source ? 9'hb6 : _GEN_183; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_185 = 9'hb7 == auto_in_a_bits_source ? 9'hb7 : _GEN_184; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_186 = 9'hb8 == auto_in_a_bits_source ? 9'hb8 : _GEN_185; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_187 = 9'hb9 == auto_in_a_bits_source ? 9'hb9 : _GEN_186; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_188 = 9'hba == auto_in_a_bits_source ? 9'hba : _GEN_187; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_189 = 9'hbb == auto_in_a_bits_source ? 9'hbb : _GEN_188; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_190 = 9'hbc == auto_in_a_bits_source ? 9'hbc : _GEN_189; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_191 = 9'hbd == auto_in_a_bits_source ? 9'hbd : _GEN_190; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_192 = 9'hbe == auto_in_a_bits_source ? 9'hbe : _GEN_191; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_193 = 9'hbf == auto_in_a_bits_source ? 9'hbf : _GEN_192; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_194 = 9'hc0 == auto_in_a_bits_source ? 9'hc0 : _GEN_193; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_195 = 9'hc1 == auto_in_a_bits_source ? 9'hc1 : _GEN_194; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_196 = 9'hc2 == auto_in_a_bits_source ? 9'hc2 : _GEN_195; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_197 = 9'hc3 == auto_in_a_bits_source ? 9'hc3 : _GEN_196; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_198 = 9'hc4 == auto_in_a_bits_source ? 9'hc4 : _GEN_197; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_199 = 9'hc5 == auto_in_a_bits_source ? 9'hc5 : _GEN_198; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_200 = 9'hc6 == auto_in_a_bits_source ? 9'hc6 : _GEN_199; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_201 = 9'hc7 == auto_in_a_bits_source ? 9'hc7 : _GEN_200; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_202 = 9'hc8 == auto_in_a_bits_source ? 9'hc8 : _GEN_201; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_203 = 9'hc9 == auto_in_a_bits_source ? 9'hc9 : _GEN_202; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_204 = 9'hca == auto_in_a_bits_source ? 9'hca : _GEN_203; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_205 = 9'hcb == auto_in_a_bits_source ? 9'hcb : _GEN_204; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_206 = 9'hcc == auto_in_a_bits_source ? 9'hcc : _GEN_205; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_207 = 9'hcd == auto_in_a_bits_source ? 9'hcd : _GEN_206; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_208 = 9'hce == auto_in_a_bits_source ? 9'hce : _GEN_207; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_209 = 9'hcf == auto_in_a_bits_source ? 9'hcf : _GEN_208; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_210 = 9'hd0 == auto_in_a_bits_source ? 9'hd0 : _GEN_209; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_211 = 9'hd1 == auto_in_a_bits_source ? 9'hd1 : _GEN_210; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_212 = 9'hd2 == auto_in_a_bits_source ? 9'hd2 : _GEN_211; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_213 = 9'hd3 == auto_in_a_bits_source ? 9'hd3 : _GEN_212; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_214 = 9'hd4 == auto_in_a_bits_source ? 9'hd4 : _GEN_213; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_215 = 9'hd5 == auto_in_a_bits_source ? 9'hd5 : _GEN_214; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_216 = 9'hd6 == auto_in_a_bits_source ? 9'hd6 : _GEN_215; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_217 = 9'hd7 == auto_in_a_bits_source ? 9'hd7 : _GEN_216; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_218 = 9'hd8 == auto_in_a_bits_source ? 9'hd8 : _GEN_217; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_219 = 9'hd9 == auto_in_a_bits_source ? 9'hd9 : _GEN_218; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_220 = 9'hda == auto_in_a_bits_source ? 9'hda : _GEN_219; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_221 = 9'hdb == auto_in_a_bits_source ? 9'hdb : _GEN_220; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_222 = 9'hdc == auto_in_a_bits_source ? 9'hdc : _GEN_221; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_223 = 9'hdd == auto_in_a_bits_source ? 9'hdd : _GEN_222; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_224 = 9'hde == auto_in_a_bits_source ? 9'hde : _GEN_223; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_225 = 9'hdf == auto_in_a_bits_source ? 9'hdf : _GEN_224; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_226 = 9'he0 == auto_in_a_bits_source ? 9'he0 : _GEN_225; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_227 = 9'he1 == auto_in_a_bits_source ? 9'he1 : _GEN_226; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_228 = 9'he2 == auto_in_a_bits_source ? 9'he2 : _GEN_227; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_229 = 9'he3 == auto_in_a_bits_source ? 9'he3 : _GEN_228; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_230 = 9'he4 == auto_in_a_bits_source ? 9'he4 : _GEN_229; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_231 = 9'he5 == auto_in_a_bits_source ? 9'he5 : _GEN_230; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_232 = 9'he6 == auto_in_a_bits_source ? 9'he6 : _GEN_231; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_233 = 9'he7 == auto_in_a_bits_source ? 9'he7 : _GEN_232; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_234 = 9'he8 == auto_in_a_bits_source ? 9'he8 : _GEN_233; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_235 = 9'he9 == auto_in_a_bits_source ? 9'he9 : _GEN_234; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_236 = 9'hea == auto_in_a_bits_source ? 9'hea : _GEN_235; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_237 = 9'heb == auto_in_a_bits_source ? 9'heb : _GEN_236; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_238 = 9'hec == auto_in_a_bits_source ? 9'hec : _GEN_237; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_239 = 9'hed == auto_in_a_bits_source ? 9'hed : _GEN_238; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_240 = 9'hee == auto_in_a_bits_source ? 9'hee : _GEN_239; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_241 = 9'hef == auto_in_a_bits_source ? 9'hef : _GEN_240; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_242 = 9'hf0 == auto_in_a_bits_source ? 9'hf0 : _GEN_241; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_243 = 9'hf1 == auto_in_a_bits_source ? 9'hf1 : _GEN_242; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_244 = 9'hf2 == auto_in_a_bits_source ? 9'hf2 : _GEN_243; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_245 = 9'hf3 == auto_in_a_bits_source ? 9'hf3 : _GEN_244; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_246 = 9'hf4 == auto_in_a_bits_source ? 9'hf4 : _GEN_245; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_247 = 9'hf5 == auto_in_a_bits_source ? 9'hf5 : _GEN_246; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_248 = 9'hf6 == auto_in_a_bits_source ? 9'hf6 : _GEN_247; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_249 = 9'hf7 == auto_in_a_bits_source ? 9'hf7 : _GEN_248; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_250 = 9'hf8 == auto_in_a_bits_source ? 9'hf8 : _GEN_249; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_251 = 9'hf9 == auto_in_a_bits_source ? 9'hf9 : _GEN_250; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_252 = 9'hfa == auto_in_a_bits_source ? 9'hfa : _GEN_251; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_253 = 9'hfb == auto_in_a_bits_source ? 9'hfb : _GEN_252; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_254 = 9'hfc == auto_in_a_bits_source ? 9'hfc : _GEN_253; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_255 = 9'hfd == auto_in_a_bits_source ? 9'hfd : _GEN_254; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_256 = 9'hfe == auto_in_a_bits_source ? 9'hfe : _GEN_255; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_257 = 9'hff == auto_in_a_bits_source ? 9'hff : _GEN_256; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_258 = 9'h100 == auto_in_a_bits_source ? 9'h100 : _GEN_257; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_259 = 9'h101 == auto_in_a_bits_source ? 9'h101 : _GEN_258; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_260 = 9'h102 == auto_in_a_bits_source ? 9'h102 : _GEN_259; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_261 = 9'h103 == auto_in_a_bits_source ? 9'h103 : _GEN_260; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_262 = 9'h104 == auto_in_a_bits_source ? 9'h104 : _GEN_261; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_263 = 9'h105 == auto_in_a_bits_source ? 9'h105 : _GEN_262; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_264 = 9'h106 == auto_in_a_bits_source ? 9'h106 : _GEN_263; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_265 = 9'h107 == auto_in_a_bits_source ? 9'h107 : _GEN_264; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_266 = 9'h108 == auto_in_a_bits_source ? 9'h108 : _GEN_265; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_267 = 9'h109 == auto_in_a_bits_source ? 9'h109 : _GEN_266; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_268 = 9'h10a == auto_in_a_bits_source ? 9'h10a : _GEN_267; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_269 = 9'h10b == auto_in_a_bits_source ? 9'h10b : _GEN_268; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_270 = 9'h10c == auto_in_a_bits_source ? 9'h10c : _GEN_269; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_271 = 9'h10d == auto_in_a_bits_source ? 9'h10d : _GEN_270; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_272 = 9'h10e == auto_in_a_bits_source ? 9'h10e : _GEN_271; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_273 = 9'h10f == auto_in_a_bits_source ? 9'h10f : _GEN_272; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_274 = 9'h110 == auto_in_a_bits_source ? 9'h110 : _GEN_273; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_275 = 9'h111 == auto_in_a_bits_source ? 9'h111 : _GEN_274; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_276 = 9'h112 == auto_in_a_bits_source ? 9'h112 : _GEN_275; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_277 = 9'h113 == auto_in_a_bits_source ? 9'h113 : _GEN_276; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_278 = 9'h114 == auto_in_a_bits_source ? 9'h114 : _GEN_277; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_279 = 9'h115 == auto_in_a_bits_source ? 9'h115 : _GEN_278; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_280 = 9'h116 == auto_in_a_bits_source ? 9'h116 : _GEN_279; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_281 = 9'h117 == auto_in_a_bits_source ? 9'h117 : _GEN_280; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_282 = 9'h118 == auto_in_a_bits_source ? 9'h118 : _GEN_281; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_283 = 9'h119 == auto_in_a_bits_source ? 9'h119 : _GEN_282; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_284 = 9'h11a == auto_in_a_bits_source ? 9'h11a : _GEN_283; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_285 = 9'h11b == auto_in_a_bits_source ? 9'h11b : _GEN_284; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_286 = 9'h11c == auto_in_a_bits_source ? 9'h11c : _GEN_285; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_287 = 9'h11d == auto_in_a_bits_source ? 9'h11d : _GEN_286; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_288 = 9'h11e == auto_in_a_bits_source ? 9'h11e : _GEN_287; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_289 = 9'h11f == auto_in_a_bits_source ? 9'h11f : _GEN_288; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_290 = 9'h120 == auto_in_a_bits_source ? 9'h120 : _GEN_289; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_291 = 9'h121 == auto_in_a_bits_source ? 9'h121 : _GEN_290; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_292 = 9'h122 == auto_in_a_bits_source ? 9'h122 : _GEN_291; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_293 = 9'h123 == auto_in_a_bits_source ? 9'h123 : _GEN_292; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_294 = 9'h124 == auto_in_a_bits_source ? 9'h124 : _GEN_293; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_295 = 9'h125 == auto_in_a_bits_source ? 9'h125 : _GEN_294; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_296 = 9'h126 == auto_in_a_bits_source ? 9'h126 : _GEN_295; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_297 = 9'h127 == auto_in_a_bits_source ? 9'h127 : _GEN_296; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_298 = 9'h128 == auto_in_a_bits_source ? 9'h128 : _GEN_297; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_299 = 9'h129 == auto_in_a_bits_source ? 9'h129 : _GEN_298; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_300 = 9'h12a == auto_in_a_bits_source ? 9'h12a : _GEN_299; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_301 = 9'h12b == auto_in_a_bits_source ? 9'h12b : _GEN_300; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_302 = 9'h12c == auto_in_a_bits_source ? 9'h12c : _GEN_301; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_303 = 9'h12d == auto_in_a_bits_source ? 9'h12d : _GEN_302; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_304 = 9'h12e == auto_in_a_bits_source ? 9'h12e : _GEN_303; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_305 = 9'h12f == auto_in_a_bits_source ? 9'h12f : _GEN_304; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_306 = 9'h130 == auto_in_a_bits_source ? 9'h130 : _GEN_305; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_307 = 9'h131 == auto_in_a_bits_source ? 9'h131 : _GEN_306; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_308 = 9'h132 == auto_in_a_bits_source ? 9'h132 : _GEN_307; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_309 = 9'h133 == auto_in_a_bits_source ? 9'h133 : _GEN_308; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_310 = 9'h134 == auto_in_a_bits_source ? 9'h134 : _GEN_309; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_311 = 9'h135 == auto_in_a_bits_source ? 9'h135 : _GEN_310; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_312 = 9'h136 == auto_in_a_bits_source ? 9'h136 : _GEN_311; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_313 = 9'h137 == auto_in_a_bits_source ? 9'h137 : _GEN_312; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_314 = 9'h138 == auto_in_a_bits_source ? 9'h138 : _GEN_313; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_315 = 9'h139 == auto_in_a_bits_source ? 9'h139 : _GEN_314; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_316 = 9'h13a == auto_in_a_bits_source ? 9'h13a : _GEN_315; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_317 = 9'h13b == auto_in_a_bits_source ? 9'h13b : _GEN_316; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_318 = 9'h13c == auto_in_a_bits_source ? 9'h13c : _GEN_317; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_319 = 9'h13d == auto_in_a_bits_source ? 9'h13d : _GEN_318; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_320 = 9'h13e == auto_in_a_bits_source ? 9'h13e : _GEN_319; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_321 = 9'h13f == auto_in_a_bits_source ? 9'h13f : _GEN_320; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_322 = 9'h140 == auto_in_a_bits_source ? 9'h140 : _GEN_321; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_323 = 9'h141 == auto_in_a_bits_source ? 9'h141 : _GEN_322; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_324 = 9'h142 == auto_in_a_bits_source ? 9'h142 : _GEN_323; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_325 = 9'h143 == auto_in_a_bits_source ? 9'h143 : _GEN_324; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_326 = 9'h144 == auto_in_a_bits_source ? 9'h144 : _GEN_325; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_327 = 9'h145 == auto_in_a_bits_source ? 9'h145 : _GEN_326; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_328 = 9'h146 == auto_in_a_bits_source ? 9'h146 : _GEN_327; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_329 = 9'h147 == auto_in_a_bits_source ? 9'h147 : _GEN_328; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_330 = 9'h148 == auto_in_a_bits_source ? 9'h148 : _GEN_329; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_331 = 9'h149 == auto_in_a_bits_source ? 9'h149 : _GEN_330; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_332 = 9'h14a == auto_in_a_bits_source ? 9'h14a : _GEN_331; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_333 = 9'h14b == auto_in_a_bits_source ? 9'h14b : _GEN_332; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_334 = 9'h14c == auto_in_a_bits_source ? 9'h14c : _GEN_333; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_335 = 9'h14d == auto_in_a_bits_source ? 9'h14d : _GEN_334; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_336 = 9'h14e == auto_in_a_bits_source ? 9'h14e : _GEN_335; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_337 = 9'h14f == auto_in_a_bits_source ? 9'h14f : _GEN_336; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_338 = 9'h150 == auto_in_a_bits_source ? 9'h150 : _GEN_337; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_339 = 9'h151 == auto_in_a_bits_source ? 9'h151 : _GEN_338; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_340 = 9'h152 == auto_in_a_bits_source ? 9'h152 : _GEN_339; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_341 = 9'h153 == auto_in_a_bits_source ? 9'h153 : _GEN_340; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_342 = 9'h154 == auto_in_a_bits_source ? 9'h154 : _GEN_341; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_343 = 9'h155 == auto_in_a_bits_source ? 9'h155 : _GEN_342; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_344 = 9'h156 == auto_in_a_bits_source ? 9'h156 : _GEN_343; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_345 = 9'h157 == auto_in_a_bits_source ? 9'h157 : _GEN_344; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_346 = 9'h158 == auto_in_a_bits_source ? 9'h158 : _GEN_345; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_347 = 9'h159 == auto_in_a_bits_source ? 9'h159 : _GEN_346; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_348 = 9'h15a == auto_in_a_bits_source ? 9'h15a : _GEN_347; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_349 = 9'h15b == auto_in_a_bits_source ? 9'h15b : _GEN_348; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_350 = 9'h15c == auto_in_a_bits_source ? 9'h15c : _GEN_349; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_351 = 9'h15d == auto_in_a_bits_source ? 9'h15d : _GEN_350; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_352 = 9'h15e == auto_in_a_bits_source ? 9'h15e : _GEN_351; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_353 = 9'h15f == auto_in_a_bits_source ? 9'h15f : _GEN_352; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_354 = 9'h160 == auto_in_a_bits_source ? 9'h160 : _GEN_353; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_355 = 9'h161 == auto_in_a_bits_source ? 9'h161 : _GEN_354; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_356 = 9'h162 == auto_in_a_bits_source ? 9'h162 : _GEN_355; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_357 = 9'h163 == auto_in_a_bits_source ? 9'h163 : _GEN_356; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_358 = 9'h164 == auto_in_a_bits_source ? 9'h164 : _GEN_357; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_359 = 9'h165 == auto_in_a_bits_source ? 9'h165 : _GEN_358; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_360 = 9'h166 == auto_in_a_bits_source ? 9'h166 : _GEN_359; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_361 = 9'h167 == auto_in_a_bits_source ? 9'h167 : _GEN_360; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_362 = 9'h168 == auto_in_a_bits_source ? 9'h168 : _GEN_361; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_363 = 9'h169 == auto_in_a_bits_source ? 9'h169 : _GEN_362; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_364 = 9'h16a == auto_in_a_bits_source ? 9'h16a : _GEN_363; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_365 = 9'h16b == auto_in_a_bits_source ? 9'h16b : _GEN_364; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_366 = 9'h16c == auto_in_a_bits_source ? 9'h16c : _GEN_365; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_367 = 9'h16d == auto_in_a_bits_source ? 9'h16d : _GEN_366; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_368 = 9'h16e == auto_in_a_bits_source ? 9'h16e : _GEN_367; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_369 = 9'h16f == auto_in_a_bits_source ? 9'h16f : _GEN_368; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_370 = 9'h170 == auto_in_a_bits_source ? 9'h170 : _GEN_369; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_371 = 9'h171 == auto_in_a_bits_source ? 9'h171 : _GEN_370; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_372 = 9'h172 == auto_in_a_bits_source ? 9'h172 : _GEN_371; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_373 = 9'h173 == auto_in_a_bits_source ? 9'h173 : _GEN_372; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_374 = 9'h174 == auto_in_a_bits_source ? 9'h174 : _GEN_373; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_375 = 9'h175 == auto_in_a_bits_source ? 9'h175 : _GEN_374; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_376 = 9'h176 == auto_in_a_bits_source ? 9'h176 : _GEN_375; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_377 = 9'h177 == auto_in_a_bits_source ? 9'h177 : _GEN_376; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_378 = 9'h178 == auto_in_a_bits_source ? 9'h178 : _GEN_377; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_379 = 9'h179 == auto_in_a_bits_source ? 9'h179 : _GEN_378; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_380 = 9'h17a == auto_in_a_bits_source ? 9'h17a : _GEN_379; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_381 = 9'h17b == auto_in_a_bits_source ? 9'h17b : _GEN_380; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_382 = 9'h17c == auto_in_a_bits_source ? 9'h17c : _GEN_381; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_383 = 9'h17d == auto_in_a_bits_source ? 9'h17d : _GEN_382; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_384 = 9'h17e == auto_in_a_bits_source ? 9'h17e : _GEN_383; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_385 = 9'h17f == auto_in_a_bits_source ? 9'h17f : _GEN_384; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_386 = 9'h180 == auto_in_a_bits_source ? 9'h180 : _GEN_385; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_387 = 9'h181 == auto_in_a_bits_source ? 9'h181 : _GEN_386; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_388 = 9'h182 == auto_in_a_bits_source ? 9'h182 : _GEN_387; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_389 = 9'h183 == auto_in_a_bits_source ? 9'h183 : _GEN_388; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_390 = 9'h184 == auto_in_a_bits_source ? 9'h184 : _GEN_389; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_391 = 9'h185 == auto_in_a_bits_source ? 9'h185 : _GEN_390; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_392 = 9'h186 == auto_in_a_bits_source ? 9'h186 : _GEN_391; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_393 = 9'h187 == auto_in_a_bits_source ? 9'h187 : _GEN_392; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_394 = 9'h188 == auto_in_a_bits_source ? 9'h188 : _GEN_393; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_395 = 9'h189 == auto_in_a_bits_source ? 9'h189 : _GEN_394; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_396 = 9'h18a == auto_in_a_bits_source ? 9'h18a : _GEN_395; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_397 = 9'h18b == auto_in_a_bits_source ? 9'h18b : _GEN_396; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_398 = 9'h18c == auto_in_a_bits_source ? 9'h18c : _GEN_397; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_399 = 9'h18d == auto_in_a_bits_source ? 9'h18d : _GEN_398; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_400 = 9'h18e == auto_in_a_bits_source ? 9'h18e : _GEN_399; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_401 = 9'h18f == auto_in_a_bits_source ? 9'h18f : _GEN_400; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_402 = 9'h190 == auto_in_a_bits_source ? 9'h190 : _GEN_401; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_403 = 9'h191 == auto_in_a_bits_source ? 9'h191 : _GEN_402; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_404 = 9'h192 == auto_in_a_bits_source ? 9'h192 : _GEN_403; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_405 = 9'h193 == auto_in_a_bits_source ? 9'h193 : _GEN_404; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_406 = 9'h194 == auto_in_a_bits_source ? 9'h194 : _GEN_405; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_407 = 9'h195 == auto_in_a_bits_source ? 9'h195 : _GEN_406; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_408 = 9'h196 == auto_in_a_bits_source ? 9'h196 : _GEN_407; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_409 = 9'h197 == auto_in_a_bits_source ? 9'h197 : _GEN_408; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_410 = 9'h198 == auto_in_a_bits_source ? 9'h198 : _GEN_409; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_411 = 9'h199 == auto_in_a_bits_source ? 9'h199 : _GEN_410; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_412 = 9'h19a == auto_in_a_bits_source ? 9'h19a : _GEN_411; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_413 = 9'h19b == auto_in_a_bits_source ? 9'h19b : _GEN_412; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_414 = 9'h19c == auto_in_a_bits_source ? 9'h19c : _GEN_413; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_415 = 9'h19d == auto_in_a_bits_source ? 9'h19d : _GEN_414; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_416 = 9'h19e == auto_in_a_bits_source ? 9'h19e : _GEN_415; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_417 = 9'h19f == auto_in_a_bits_source ? 9'h19f : _GEN_416; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_418 = 9'h1a0 == auto_in_a_bits_source ? 9'h1a0 : _GEN_417; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_419 = 9'h1a1 == auto_in_a_bits_source ? 9'h1a1 : _GEN_418; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_420 = 9'h1a2 == auto_in_a_bits_source ? 9'h1a2 : _GEN_419; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_421 = 9'h1a3 == auto_in_a_bits_source ? 9'h1a3 : _GEN_420; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_422 = 9'h1a4 == auto_in_a_bits_source ? 9'h1a4 : _GEN_421; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_423 = 9'h1a5 == auto_in_a_bits_source ? 9'h1a5 : _GEN_422; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_424 = 9'h1a6 == auto_in_a_bits_source ? 9'h1a6 : _GEN_423; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_425 = 9'h1a7 == auto_in_a_bits_source ? 9'h1a7 : _GEN_424; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_426 = 9'h1a8 == auto_in_a_bits_source ? 9'h1a8 : _GEN_425; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_427 = 9'h1a9 == auto_in_a_bits_source ? 9'h1a9 : _GEN_426; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_428 = 9'h1aa == auto_in_a_bits_source ? 9'h1aa : _GEN_427; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_429 = 9'h1ab == auto_in_a_bits_source ? 9'h1ab : _GEN_428; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_430 = 9'h1ac == auto_in_a_bits_source ? 9'h1ac : _GEN_429; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_431 = 9'h1ad == auto_in_a_bits_source ? 9'h1ad : _GEN_430; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_432 = 9'h1ae == auto_in_a_bits_source ? 9'h1ae : _GEN_431; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_433 = 9'h1af == auto_in_a_bits_source ? 9'h1af : _GEN_432; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_434 = 9'h1b0 == auto_in_a_bits_source ? 9'h1b0 : _GEN_433; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_435 = 9'h1b1 == auto_in_a_bits_source ? 9'h1b1 : _GEN_434; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_436 = 9'h1b2 == auto_in_a_bits_source ? 9'h1b2 : _GEN_435; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_437 = 9'h1b3 == auto_in_a_bits_source ? 9'h1b3 : _GEN_436; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_438 = 9'h1b4 == auto_in_a_bits_source ? 9'h1b4 : _GEN_437; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_439 = 9'h1b5 == auto_in_a_bits_source ? 9'h1b5 : _GEN_438; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_440 = 9'h1b6 == auto_in_a_bits_source ? 9'h1b6 : _GEN_439; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_441 = 9'h1b7 == auto_in_a_bits_source ? 9'h1b7 : _GEN_440; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_442 = 9'h1b8 == auto_in_a_bits_source ? 9'h1b8 : _GEN_441; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_443 = 9'h1b9 == auto_in_a_bits_source ? 9'h1b9 : _GEN_442; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_444 = 9'h1ba == auto_in_a_bits_source ? 9'h1ba : _GEN_443; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_445 = 9'h1bb == auto_in_a_bits_source ? 9'h1bb : _GEN_444; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_446 = 9'h1bc == auto_in_a_bits_source ? 9'h1bc : _GEN_445; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_447 = 9'h1bd == auto_in_a_bits_source ? 9'h1bd : _GEN_446; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_448 = 9'h1be == auto_in_a_bits_source ? 9'h1be : _GEN_447; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_449 = 9'h1bf == auto_in_a_bits_source ? 9'h1bf : _GEN_448; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_450 = 9'h1c0 == auto_in_a_bits_source ? 9'h1c0 : _GEN_449; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_451 = 9'h1c1 == auto_in_a_bits_source ? 9'h1c1 : _GEN_450; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_452 = 9'h1c2 == auto_in_a_bits_source ? 9'h1c2 : _GEN_451; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_453 = 9'h1c3 == auto_in_a_bits_source ? 9'h1c3 : _GEN_452; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_454 = 9'h1c4 == auto_in_a_bits_source ? 9'h1c4 : _GEN_453; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_455 = 9'h1c5 == auto_in_a_bits_source ? 9'h1c5 : _GEN_454; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_456 = 9'h1c6 == auto_in_a_bits_source ? 9'h1c6 : _GEN_455; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_457 = 9'h1c7 == auto_in_a_bits_source ? 9'h1c7 : _GEN_456; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_458 = 9'h1c8 == auto_in_a_bits_source ? 9'h1c8 : _GEN_457; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_459 = 9'h1c9 == auto_in_a_bits_source ? 9'h1c9 : _GEN_458; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_460 = 9'h1ca == auto_in_a_bits_source ? 9'h1ca : _GEN_459; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_461 = 9'h1cb == auto_in_a_bits_source ? 9'h1cb : _GEN_460; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_462 = 9'h1cc == auto_in_a_bits_source ? 9'h1cc : _GEN_461; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_463 = 9'h1cd == auto_in_a_bits_source ? 9'h1cd : _GEN_462; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_464 = 9'h1ce == auto_in_a_bits_source ? 9'h1ce : _GEN_463; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_465 = 9'h1cf == auto_in_a_bits_source ? 9'h1cf : _GEN_464; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_466 = 9'h1d0 == auto_in_a_bits_source ? 9'h1d0 : _GEN_465; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_467 = 9'h1d1 == auto_in_a_bits_source ? 9'h1d1 : _GEN_466; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_468 = 9'h1d2 == auto_in_a_bits_source ? 9'h1d2 : _GEN_467; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_469 = 9'h1d3 == auto_in_a_bits_source ? 9'h1d3 : _GEN_468; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_470 = 9'h1d4 == auto_in_a_bits_source ? 9'h1d4 : _GEN_469; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_471 = 9'h1d5 == auto_in_a_bits_source ? 9'h1d5 : _GEN_470; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_472 = 9'h1d6 == auto_in_a_bits_source ? 9'h1d6 : _GEN_471; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_473 = 9'h1d7 == auto_in_a_bits_source ? 9'h1d7 : _GEN_472; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_474 = 9'h1d8 == auto_in_a_bits_source ? 9'h1d8 : _GEN_473; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_475 = 9'h1d9 == auto_in_a_bits_source ? 9'h1d9 : _GEN_474; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_476 = 9'h1da == auto_in_a_bits_source ? 9'h1da : _GEN_475; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_477 = 9'h1db == auto_in_a_bits_source ? 9'h1db : _GEN_476; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_478 = 9'h1dc == auto_in_a_bits_source ? 9'h1dc : _GEN_477; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_479 = 9'h1dd == auto_in_a_bits_source ? 9'h1dd : _GEN_478; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_480 = 9'h1de == auto_in_a_bits_source ? 9'h1de : _GEN_479; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_481 = 9'h1df == auto_in_a_bits_source ? 9'h1df : _GEN_480; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_482 = 9'h1e0 == auto_in_a_bits_source ? 9'h1e0 : _GEN_481; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_483 = 9'h1e1 == auto_in_a_bits_source ? 9'h1e1 : _GEN_482; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_484 = 9'h1e2 == auto_in_a_bits_source ? 9'h1e2 : _GEN_483; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_485 = 9'h1e3 == auto_in_a_bits_source ? 9'h1e3 : _GEN_484; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_486 = 9'h1e4 == auto_in_a_bits_source ? 9'h1e4 : _GEN_485; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_487 = 9'h1e5 == auto_in_a_bits_source ? 9'h1e5 : _GEN_486; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_488 = 9'h1e6 == auto_in_a_bits_source ? 9'h1e6 : _GEN_487; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_489 = 9'h1e7 == auto_in_a_bits_source ? 9'h1e7 : _GEN_488; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_490 = 9'h1e8 == auto_in_a_bits_source ? 9'h1e8 : _GEN_489; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_491 = 9'h1e9 == auto_in_a_bits_source ? 9'h1e9 : _GEN_490; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_492 = 9'h1ea == auto_in_a_bits_source ? 9'h1ea : _GEN_491; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_493 = 9'h1eb == auto_in_a_bits_source ? 9'h1eb : _GEN_492; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_494 = 9'h1ec == auto_in_a_bits_source ? 9'h1ec : _GEN_493; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_495 = 9'h1ed == auto_in_a_bits_source ? 9'h1ed : _GEN_494; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_496 = 9'h1ee == auto_in_a_bits_source ? 9'h1ee : _GEN_495; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_497 = 9'h1ef == auto_in_a_bits_source ? 9'h1ef : _GEN_496; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_498 = 9'h1f0 == auto_in_a_bits_source ? 9'h1f0 : _GEN_497; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_499 = 9'h1f1 == auto_in_a_bits_source ? 9'h1f1 : _GEN_498; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_500 = 9'h1f2 == auto_in_a_bits_source ? 9'h1f2 : _GEN_499; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_501 = 9'h1f3 == auto_in_a_bits_source ? 9'h1f3 : _GEN_500; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_502 = 9'h1f4 == auto_in_a_bits_source ? 9'h1f4 : _GEN_501; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_503 = 9'h1f5 == auto_in_a_bits_source ? 9'h1f5 : _GEN_502; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_504 = 9'h1f6 == auto_in_a_bits_source ? 9'h1f6 : _GEN_503; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_505 = 9'h1f7 == auto_in_a_bits_source ? 9'h1f7 : _GEN_504; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_506 = 9'h1f8 == auto_in_a_bits_source ? 9'h1f8 : _GEN_505; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_507 = 9'h1f9 == auto_in_a_bits_source ? 9'h1f9 : _GEN_506; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_508 = 9'h1fa == auto_in_a_bits_source ? 9'h1fa : _GEN_507; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_509 = 9'h1fb == auto_in_a_bits_source ? 9'h1fb : _GEN_508; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_510 = 9'h1fc == auto_in_a_bits_source ? 9'h1fc : _GEN_509; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_511 = 9'h1fd == auto_in_a_bits_source ? 9'h1fd : _GEN_510; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] _GEN_512 = 9'h1fe == auto_in_a_bits_source ? 9'h1fe : _GEN_511; // @[ToAXI4.scala 166:{17,17}]
  wire [8:0] out_arw_bits_id = 9'h1ff == auto_in_a_bits_source ? 9'h1ff : _GEN_512; // @[ToAXI4.scala 166:{17,17}]
  wire [17:0] _out_arw_bits_len_T_1 = 18'h7ff << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [10:0] _out_arw_bits_len_T_3 = ~_out_arw_bits_len_T_1[10:0]; // @[package.scala 234:46]
  wire  prot_1 = ~auto_in_a_bits_user_amba_prot_secure; // @[ToAXI4.scala 185:20]
  wire [1:0] out_arw_bits_prot_hi = {auto_in_a_bits_user_amba_prot_fetch,prot_1}; // @[Cat.scala 31:58]
  wire [1:0] out_arw_bits_cache_lo = {auto_in_a_bits_user_amba_prot_modifiable,auto_in_a_bits_user_amba_prot_bufferable}
    ; // @[Cat.scala 31:58]
  wire [1:0] out_arw_bits_cache_hi = {auto_in_a_bits_user_amba_prot_writealloc,auto_in_a_bits_user_amba_prot_readalloc}; // @[Cat.scala 31:58]
  wire  _out_arw_valid_T_1 = _bundleIn_0_a_ready_T & auto_in_a_valid; // @[ToAXI4.scala 197:31]
  wire  _out_arw_valid_T_4 = a_isPut ? ~doneAW & out_w_ready : 1'h1; // @[ToAXI4.scala 197:51]
  wire  out_arw_valid = _bundleIn_0_a_ready_T & auto_in_a_valid & _out_arw_valid_T_4; // @[ToAXI4.scala 197:45]
  reg  r_holds_d; // @[ToAXI4.scala 206:30]
  reg [2:0] b_delay; // @[ToAXI4.scala 209:24]
  wire  r_wins = auto_out_r_valid & b_delay != 3'h7 | r_holds_d; // @[ToAXI4.scala 215:57]
  wire  bundleOut_0_r_ready = auto_in_d_ready & r_wins; // @[ToAXI4.scala 217:33]
  wire  _T_2 = bundleOut_0_r_ready & auto_out_r_valid; // @[Decoupled.scala 50:35]
  wire  bundleOut_0_b_ready = auto_in_d_ready & ~r_wins; // @[ToAXI4.scala 218:33]
  wire [2:0] _b_delay_T_1 = b_delay + 3'h1; // @[ToAXI4.scala 211:28]
  wire  bundleIn_0_d_valid = r_wins ? auto_out_r_valid : auto_out_b_valid; // @[ToAXI4.scala 219:24]
  reg  r_first; // @[ToAXI4.scala 224:28]
  wire  _GEN_1028 = _T_2 ? auto_out_r_bits_last : r_first; // @[ToAXI4.scala 225:27 224:28 225:37]
  wire  _r_denied_T = auto_out_r_bits_resp == 2'h3; // @[ToAXI4.scala 226:39]
  reg  r_denied_r; // @[Reg.scala 16:16]
  wire  _GEN_1029 = r_first ? _r_denied_T : r_denied_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  r_corrupt = auto_out_r_bits_resp != 2'h0; // @[ToAXI4.scala 227:39]
  wire  b_denied = auto_out_b_bits_resp != 2'h0; // @[ToAXI4.scala 228:39]
  wire  r_d_corrupt = r_corrupt | _GEN_1029; // @[ToAXI4.scala 230:100]
  wire [2:0] r_d_size = auto_out_r_bits_echo_tl_state_size[2:0]; // @[Edges.scala 771:17 774:15]
  wire [2:0] b_d_size = auto_out_b_bits_echo_tl_state_size[2:0]; // @[Edges.scala 755:17 758:15]
  wire [511:0] _a_sel_T = 512'h1 << out_arw_bits_id; // @[OneHot.scala 64:12]
  wire  a_sel_0 = _a_sel_T[0]; // @[ToAXI4.scala 242:58]
  wire  a_sel_1 = _a_sel_T[1]; // @[ToAXI4.scala 242:58]
  wire  a_sel_2 = _a_sel_T[2]; // @[ToAXI4.scala 242:58]
  wire  a_sel_3 = _a_sel_T[3]; // @[ToAXI4.scala 242:58]
  wire  a_sel_4 = _a_sel_T[4]; // @[ToAXI4.scala 242:58]
  wire  a_sel_5 = _a_sel_T[5]; // @[ToAXI4.scala 242:58]
  wire  a_sel_6 = _a_sel_T[6]; // @[ToAXI4.scala 242:58]
  wire  a_sel_7 = _a_sel_T[7]; // @[ToAXI4.scala 242:58]
  wire  a_sel_8 = _a_sel_T[8]; // @[ToAXI4.scala 242:58]
  wire  a_sel_9 = _a_sel_T[9]; // @[ToAXI4.scala 242:58]
  wire  a_sel_10 = _a_sel_T[10]; // @[ToAXI4.scala 242:58]
  wire  a_sel_11 = _a_sel_T[11]; // @[ToAXI4.scala 242:58]
  wire  a_sel_12 = _a_sel_T[12]; // @[ToAXI4.scala 242:58]
  wire  a_sel_13 = _a_sel_T[13]; // @[ToAXI4.scala 242:58]
  wire  a_sel_14 = _a_sel_T[14]; // @[ToAXI4.scala 242:58]
  wire  a_sel_15 = _a_sel_T[15]; // @[ToAXI4.scala 242:58]
  wire  a_sel_16 = _a_sel_T[16]; // @[ToAXI4.scala 242:58]
  wire  a_sel_17 = _a_sel_T[17]; // @[ToAXI4.scala 242:58]
  wire  a_sel_18 = _a_sel_T[18]; // @[ToAXI4.scala 242:58]
  wire  a_sel_19 = _a_sel_T[19]; // @[ToAXI4.scala 242:58]
  wire  a_sel_20 = _a_sel_T[20]; // @[ToAXI4.scala 242:58]
  wire  a_sel_21 = _a_sel_T[21]; // @[ToAXI4.scala 242:58]
  wire  a_sel_22 = _a_sel_T[22]; // @[ToAXI4.scala 242:58]
  wire  a_sel_23 = _a_sel_T[23]; // @[ToAXI4.scala 242:58]
  wire  a_sel_24 = _a_sel_T[24]; // @[ToAXI4.scala 242:58]
  wire  a_sel_25 = _a_sel_T[25]; // @[ToAXI4.scala 242:58]
  wire  a_sel_26 = _a_sel_T[26]; // @[ToAXI4.scala 242:58]
  wire  a_sel_27 = _a_sel_T[27]; // @[ToAXI4.scala 242:58]
  wire  a_sel_28 = _a_sel_T[28]; // @[ToAXI4.scala 242:58]
  wire  a_sel_29 = _a_sel_T[29]; // @[ToAXI4.scala 242:58]
  wire  a_sel_30 = _a_sel_T[30]; // @[ToAXI4.scala 242:58]
  wire  a_sel_31 = _a_sel_T[31]; // @[ToAXI4.scala 242:58]
  wire  a_sel_32 = _a_sel_T[32]; // @[ToAXI4.scala 242:58]
  wire  a_sel_33 = _a_sel_T[33]; // @[ToAXI4.scala 242:58]
  wire  a_sel_34 = _a_sel_T[34]; // @[ToAXI4.scala 242:58]
  wire  a_sel_35 = _a_sel_T[35]; // @[ToAXI4.scala 242:58]
  wire  a_sel_36 = _a_sel_T[36]; // @[ToAXI4.scala 242:58]
  wire  a_sel_37 = _a_sel_T[37]; // @[ToAXI4.scala 242:58]
  wire  a_sel_38 = _a_sel_T[38]; // @[ToAXI4.scala 242:58]
  wire  a_sel_39 = _a_sel_T[39]; // @[ToAXI4.scala 242:58]
  wire  a_sel_40 = _a_sel_T[40]; // @[ToAXI4.scala 242:58]
  wire  a_sel_41 = _a_sel_T[41]; // @[ToAXI4.scala 242:58]
  wire  a_sel_42 = _a_sel_T[42]; // @[ToAXI4.scala 242:58]
  wire  a_sel_43 = _a_sel_T[43]; // @[ToAXI4.scala 242:58]
  wire  a_sel_44 = _a_sel_T[44]; // @[ToAXI4.scala 242:58]
  wire  a_sel_45 = _a_sel_T[45]; // @[ToAXI4.scala 242:58]
  wire  a_sel_46 = _a_sel_T[46]; // @[ToAXI4.scala 242:58]
  wire  a_sel_47 = _a_sel_T[47]; // @[ToAXI4.scala 242:58]
  wire  a_sel_48 = _a_sel_T[48]; // @[ToAXI4.scala 242:58]
  wire  a_sel_49 = _a_sel_T[49]; // @[ToAXI4.scala 242:58]
  wire  a_sel_50 = _a_sel_T[50]; // @[ToAXI4.scala 242:58]
  wire  a_sel_51 = _a_sel_T[51]; // @[ToAXI4.scala 242:58]
  wire  a_sel_52 = _a_sel_T[52]; // @[ToAXI4.scala 242:58]
  wire  a_sel_53 = _a_sel_T[53]; // @[ToAXI4.scala 242:58]
  wire  a_sel_54 = _a_sel_T[54]; // @[ToAXI4.scala 242:58]
  wire  a_sel_55 = _a_sel_T[55]; // @[ToAXI4.scala 242:58]
  wire  a_sel_56 = _a_sel_T[56]; // @[ToAXI4.scala 242:58]
  wire  a_sel_57 = _a_sel_T[57]; // @[ToAXI4.scala 242:58]
  wire  a_sel_58 = _a_sel_T[58]; // @[ToAXI4.scala 242:58]
  wire  a_sel_59 = _a_sel_T[59]; // @[ToAXI4.scala 242:58]
  wire  a_sel_60 = _a_sel_T[60]; // @[ToAXI4.scala 242:58]
  wire  a_sel_61 = _a_sel_T[61]; // @[ToAXI4.scala 242:58]
  wire  a_sel_62 = _a_sel_T[62]; // @[ToAXI4.scala 242:58]
  wire  a_sel_63 = _a_sel_T[63]; // @[ToAXI4.scala 242:58]
  wire  a_sel_64 = _a_sel_T[64]; // @[ToAXI4.scala 242:58]
  wire  a_sel_65 = _a_sel_T[65]; // @[ToAXI4.scala 242:58]
  wire  a_sel_66 = _a_sel_T[66]; // @[ToAXI4.scala 242:58]
  wire  a_sel_67 = _a_sel_T[67]; // @[ToAXI4.scala 242:58]
  wire  a_sel_68 = _a_sel_T[68]; // @[ToAXI4.scala 242:58]
  wire  a_sel_69 = _a_sel_T[69]; // @[ToAXI4.scala 242:58]
  wire  a_sel_70 = _a_sel_T[70]; // @[ToAXI4.scala 242:58]
  wire  a_sel_71 = _a_sel_T[71]; // @[ToAXI4.scala 242:58]
  wire  a_sel_72 = _a_sel_T[72]; // @[ToAXI4.scala 242:58]
  wire  a_sel_73 = _a_sel_T[73]; // @[ToAXI4.scala 242:58]
  wire  a_sel_74 = _a_sel_T[74]; // @[ToAXI4.scala 242:58]
  wire  a_sel_75 = _a_sel_T[75]; // @[ToAXI4.scala 242:58]
  wire  a_sel_76 = _a_sel_T[76]; // @[ToAXI4.scala 242:58]
  wire  a_sel_77 = _a_sel_T[77]; // @[ToAXI4.scala 242:58]
  wire  a_sel_78 = _a_sel_T[78]; // @[ToAXI4.scala 242:58]
  wire  a_sel_79 = _a_sel_T[79]; // @[ToAXI4.scala 242:58]
  wire  a_sel_80 = _a_sel_T[80]; // @[ToAXI4.scala 242:58]
  wire  a_sel_81 = _a_sel_T[81]; // @[ToAXI4.scala 242:58]
  wire  a_sel_82 = _a_sel_T[82]; // @[ToAXI4.scala 242:58]
  wire  a_sel_83 = _a_sel_T[83]; // @[ToAXI4.scala 242:58]
  wire  a_sel_84 = _a_sel_T[84]; // @[ToAXI4.scala 242:58]
  wire  a_sel_85 = _a_sel_T[85]; // @[ToAXI4.scala 242:58]
  wire  a_sel_86 = _a_sel_T[86]; // @[ToAXI4.scala 242:58]
  wire  a_sel_87 = _a_sel_T[87]; // @[ToAXI4.scala 242:58]
  wire  a_sel_88 = _a_sel_T[88]; // @[ToAXI4.scala 242:58]
  wire  a_sel_89 = _a_sel_T[89]; // @[ToAXI4.scala 242:58]
  wire  a_sel_90 = _a_sel_T[90]; // @[ToAXI4.scala 242:58]
  wire  a_sel_91 = _a_sel_T[91]; // @[ToAXI4.scala 242:58]
  wire  a_sel_92 = _a_sel_T[92]; // @[ToAXI4.scala 242:58]
  wire  a_sel_93 = _a_sel_T[93]; // @[ToAXI4.scala 242:58]
  wire  a_sel_94 = _a_sel_T[94]; // @[ToAXI4.scala 242:58]
  wire  a_sel_95 = _a_sel_T[95]; // @[ToAXI4.scala 242:58]
  wire  a_sel_96 = _a_sel_T[96]; // @[ToAXI4.scala 242:58]
  wire  a_sel_97 = _a_sel_T[97]; // @[ToAXI4.scala 242:58]
  wire  a_sel_98 = _a_sel_T[98]; // @[ToAXI4.scala 242:58]
  wire  a_sel_99 = _a_sel_T[99]; // @[ToAXI4.scala 242:58]
  wire  a_sel_100 = _a_sel_T[100]; // @[ToAXI4.scala 242:58]
  wire  a_sel_101 = _a_sel_T[101]; // @[ToAXI4.scala 242:58]
  wire  a_sel_102 = _a_sel_T[102]; // @[ToAXI4.scala 242:58]
  wire  a_sel_103 = _a_sel_T[103]; // @[ToAXI4.scala 242:58]
  wire  a_sel_104 = _a_sel_T[104]; // @[ToAXI4.scala 242:58]
  wire  a_sel_105 = _a_sel_T[105]; // @[ToAXI4.scala 242:58]
  wire  a_sel_106 = _a_sel_T[106]; // @[ToAXI4.scala 242:58]
  wire  a_sel_107 = _a_sel_T[107]; // @[ToAXI4.scala 242:58]
  wire  a_sel_108 = _a_sel_T[108]; // @[ToAXI4.scala 242:58]
  wire  a_sel_109 = _a_sel_T[109]; // @[ToAXI4.scala 242:58]
  wire  a_sel_110 = _a_sel_T[110]; // @[ToAXI4.scala 242:58]
  wire  a_sel_111 = _a_sel_T[111]; // @[ToAXI4.scala 242:58]
  wire  a_sel_112 = _a_sel_T[112]; // @[ToAXI4.scala 242:58]
  wire  a_sel_113 = _a_sel_T[113]; // @[ToAXI4.scala 242:58]
  wire  a_sel_114 = _a_sel_T[114]; // @[ToAXI4.scala 242:58]
  wire  a_sel_115 = _a_sel_T[115]; // @[ToAXI4.scala 242:58]
  wire  a_sel_116 = _a_sel_T[116]; // @[ToAXI4.scala 242:58]
  wire  a_sel_117 = _a_sel_T[117]; // @[ToAXI4.scala 242:58]
  wire  a_sel_118 = _a_sel_T[118]; // @[ToAXI4.scala 242:58]
  wire  a_sel_119 = _a_sel_T[119]; // @[ToAXI4.scala 242:58]
  wire  a_sel_120 = _a_sel_T[120]; // @[ToAXI4.scala 242:58]
  wire  a_sel_121 = _a_sel_T[121]; // @[ToAXI4.scala 242:58]
  wire  a_sel_122 = _a_sel_T[122]; // @[ToAXI4.scala 242:58]
  wire  a_sel_123 = _a_sel_T[123]; // @[ToAXI4.scala 242:58]
  wire  a_sel_124 = _a_sel_T[124]; // @[ToAXI4.scala 242:58]
  wire  a_sel_125 = _a_sel_T[125]; // @[ToAXI4.scala 242:58]
  wire  a_sel_126 = _a_sel_T[126]; // @[ToAXI4.scala 242:58]
  wire  a_sel_127 = _a_sel_T[127]; // @[ToAXI4.scala 242:58]
  wire  a_sel_128 = _a_sel_T[128]; // @[ToAXI4.scala 242:58]
  wire  a_sel_129 = _a_sel_T[129]; // @[ToAXI4.scala 242:58]
  wire  a_sel_130 = _a_sel_T[130]; // @[ToAXI4.scala 242:58]
  wire  a_sel_131 = _a_sel_T[131]; // @[ToAXI4.scala 242:58]
  wire  a_sel_132 = _a_sel_T[132]; // @[ToAXI4.scala 242:58]
  wire  a_sel_133 = _a_sel_T[133]; // @[ToAXI4.scala 242:58]
  wire  a_sel_134 = _a_sel_T[134]; // @[ToAXI4.scala 242:58]
  wire  a_sel_135 = _a_sel_T[135]; // @[ToAXI4.scala 242:58]
  wire  a_sel_136 = _a_sel_T[136]; // @[ToAXI4.scala 242:58]
  wire  a_sel_137 = _a_sel_T[137]; // @[ToAXI4.scala 242:58]
  wire  a_sel_138 = _a_sel_T[138]; // @[ToAXI4.scala 242:58]
  wire  a_sel_139 = _a_sel_T[139]; // @[ToAXI4.scala 242:58]
  wire  a_sel_140 = _a_sel_T[140]; // @[ToAXI4.scala 242:58]
  wire  a_sel_141 = _a_sel_T[141]; // @[ToAXI4.scala 242:58]
  wire  a_sel_142 = _a_sel_T[142]; // @[ToAXI4.scala 242:58]
  wire  a_sel_143 = _a_sel_T[143]; // @[ToAXI4.scala 242:58]
  wire  a_sel_144 = _a_sel_T[144]; // @[ToAXI4.scala 242:58]
  wire  a_sel_145 = _a_sel_T[145]; // @[ToAXI4.scala 242:58]
  wire  a_sel_146 = _a_sel_T[146]; // @[ToAXI4.scala 242:58]
  wire  a_sel_147 = _a_sel_T[147]; // @[ToAXI4.scala 242:58]
  wire  a_sel_148 = _a_sel_T[148]; // @[ToAXI4.scala 242:58]
  wire  a_sel_149 = _a_sel_T[149]; // @[ToAXI4.scala 242:58]
  wire  a_sel_150 = _a_sel_T[150]; // @[ToAXI4.scala 242:58]
  wire  a_sel_151 = _a_sel_T[151]; // @[ToAXI4.scala 242:58]
  wire  a_sel_152 = _a_sel_T[152]; // @[ToAXI4.scala 242:58]
  wire  a_sel_153 = _a_sel_T[153]; // @[ToAXI4.scala 242:58]
  wire  a_sel_154 = _a_sel_T[154]; // @[ToAXI4.scala 242:58]
  wire  a_sel_155 = _a_sel_T[155]; // @[ToAXI4.scala 242:58]
  wire  a_sel_156 = _a_sel_T[156]; // @[ToAXI4.scala 242:58]
  wire  a_sel_157 = _a_sel_T[157]; // @[ToAXI4.scala 242:58]
  wire  a_sel_158 = _a_sel_T[158]; // @[ToAXI4.scala 242:58]
  wire  a_sel_159 = _a_sel_T[159]; // @[ToAXI4.scala 242:58]
  wire  a_sel_160 = _a_sel_T[160]; // @[ToAXI4.scala 242:58]
  wire  a_sel_161 = _a_sel_T[161]; // @[ToAXI4.scala 242:58]
  wire  a_sel_162 = _a_sel_T[162]; // @[ToAXI4.scala 242:58]
  wire  a_sel_163 = _a_sel_T[163]; // @[ToAXI4.scala 242:58]
  wire  a_sel_164 = _a_sel_T[164]; // @[ToAXI4.scala 242:58]
  wire  a_sel_165 = _a_sel_T[165]; // @[ToAXI4.scala 242:58]
  wire  a_sel_166 = _a_sel_T[166]; // @[ToAXI4.scala 242:58]
  wire  a_sel_167 = _a_sel_T[167]; // @[ToAXI4.scala 242:58]
  wire  a_sel_168 = _a_sel_T[168]; // @[ToAXI4.scala 242:58]
  wire  a_sel_169 = _a_sel_T[169]; // @[ToAXI4.scala 242:58]
  wire  a_sel_170 = _a_sel_T[170]; // @[ToAXI4.scala 242:58]
  wire  a_sel_171 = _a_sel_T[171]; // @[ToAXI4.scala 242:58]
  wire  a_sel_172 = _a_sel_T[172]; // @[ToAXI4.scala 242:58]
  wire  a_sel_173 = _a_sel_T[173]; // @[ToAXI4.scala 242:58]
  wire  a_sel_174 = _a_sel_T[174]; // @[ToAXI4.scala 242:58]
  wire  a_sel_175 = _a_sel_T[175]; // @[ToAXI4.scala 242:58]
  wire  a_sel_176 = _a_sel_T[176]; // @[ToAXI4.scala 242:58]
  wire  a_sel_177 = _a_sel_T[177]; // @[ToAXI4.scala 242:58]
  wire  a_sel_178 = _a_sel_T[178]; // @[ToAXI4.scala 242:58]
  wire  a_sel_179 = _a_sel_T[179]; // @[ToAXI4.scala 242:58]
  wire  a_sel_180 = _a_sel_T[180]; // @[ToAXI4.scala 242:58]
  wire  a_sel_181 = _a_sel_T[181]; // @[ToAXI4.scala 242:58]
  wire  a_sel_182 = _a_sel_T[182]; // @[ToAXI4.scala 242:58]
  wire  a_sel_183 = _a_sel_T[183]; // @[ToAXI4.scala 242:58]
  wire  a_sel_184 = _a_sel_T[184]; // @[ToAXI4.scala 242:58]
  wire  a_sel_185 = _a_sel_T[185]; // @[ToAXI4.scala 242:58]
  wire  a_sel_186 = _a_sel_T[186]; // @[ToAXI4.scala 242:58]
  wire  a_sel_187 = _a_sel_T[187]; // @[ToAXI4.scala 242:58]
  wire  a_sel_188 = _a_sel_T[188]; // @[ToAXI4.scala 242:58]
  wire  a_sel_189 = _a_sel_T[189]; // @[ToAXI4.scala 242:58]
  wire  a_sel_190 = _a_sel_T[190]; // @[ToAXI4.scala 242:58]
  wire  a_sel_191 = _a_sel_T[191]; // @[ToAXI4.scala 242:58]
  wire  a_sel_192 = _a_sel_T[192]; // @[ToAXI4.scala 242:58]
  wire  a_sel_193 = _a_sel_T[193]; // @[ToAXI4.scala 242:58]
  wire  a_sel_194 = _a_sel_T[194]; // @[ToAXI4.scala 242:58]
  wire  a_sel_195 = _a_sel_T[195]; // @[ToAXI4.scala 242:58]
  wire  a_sel_196 = _a_sel_T[196]; // @[ToAXI4.scala 242:58]
  wire  a_sel_197 = _a_sel_T[197]; // @[ToAXI4.scala 242:58]
  wire  a_sel_198 = _a_sel_T[198]; // @[ToAXI4.scala 242:58]
  wire  a_sel_199 = _a_sel_T[199]; // @[ToAXI4.scala 242:58]
  wire  a_sel_200 = _a_sel_T[200]; // @[ToAXI4.scala 242:58]
  wire  a_sel_201 = _a_sel_T[201]; // @[ToAXI4.scala 242:58]
  wire  a_sel_202 = _a_sel_T[202]; // @[ToAXI4.scala 242:58]
  wire  a_sel_203 = _a_sel_T[203]; // @[ToAXI4.scala 242:58]
  wire  a_sel_204 = _a_sel_T[204]; // @[ToAXI4.scala 242:58]
  wire  a_sel_205 = _a_sel_T[205]; // @[ToAXI4.scala 242:58]
  wire  a_sel_206 = _a_sel_T[206]; // @[ToAXI4.scala 242:58]
  wire  a_sel_207 = _a_sel_T[207]; // @[ToAXI4.scala 242:58]
  wire  a_sel_208 = _a_sel_T[208]; // @[ToAXI4.scala 242:58]
  wire  a_sel_209 = _a_sel_T[209]; // @[ToAXI4.scala 242:58]
  wire  a_sel_210 = _a_sel_T[210]; // @[ToAXI4.scala 242:58]
  wire  a_sel_211 = _a_sel_T[211]; // @[ToAXI4.scala 242:58]
  wire  a_sel_212 = _a_sel_T[212]; // @[ToAXI4.scala 242:58]
  wire  a_sel_213 = _a_sel_T[213]; // @[ToAXI4.scala 242:58]
  wire  a_sel_214 = _a_sel_T[214]; // @[ToAXI4.scala 242:58]
  wire  a_sel_215 = _a_sel_T[215]; // @[ToAXI4.scala 242:58]
  wire  a_sel_216 = _a_sel_T[216]; // @[ToAXI4.scala 242:58]
  wire  a_sel_217 = _a_sel_T[217]; // @[ToAXI4.scala 242:58]
  wire  a_sel_218 = _a_sel_T[218]; // @[ToAXI4.scala 242:58]
  wire  a_sel_219 = _a_sel_T[219]; // @[ToAXI4.scala 242:58]
  wire  a_sel_220 = _a_sel_T[220]; // @[ToAXI4.scala 242:58]
  wire  a_sel_221 = _a_sel_T[221]; // @[ToAXI4.scala 242:58]
  wire  a_sel_222 = _a_sel_T[222]; // @[ToAXI4.scala 242:58]
  wire  a_sel_223 = _a_sel_T[223]; // @[ToAXI4.scala 242:58]
  wire  a_sel_224 = _a_sel_T[224]; // @[ToAXI4.scala 242:58]
  wire  a_sel_225 = _a_sel_T[225]; // @[ToAXI4.scala 242:58]
  wire  a_sel_226 = _a_sel_T[226]; // @[ToAXI4.scala 242:58]
  wire  a_sel_227 = _a_sel_T[227]; // @[ToAXI4.scala 242:58]
  wire  a_sel_228 = _a_sel_T[228]; // @[ToAXI4.scala 242:58]
  wire  a_sel_229 = _a_sel_T[229]; // @[ToAXI4.scala 242:58]
  wire  a_sel_230 = _a_sel_T[230]; // @[ToAXI4.scala 242:58]
  wire  a_sel_231 = _a_sel_T[231]; // @[ToAXI4.scala 242:58]
  wire  a_sel_232 = _a_sel_T[232]; // @[ToAXI4.scala 242:58]
  wire  a_sel_233 = _a_sel_T[233]; // @[ToAXI4.scala 242:58]
  wire  a_sel_234 = _a_sel_T[234]; // @[ToAXI4.scala 242:58]
  wire  a_sel_235 = _a_sel_T[235]; // @[ToAXI4.scala 242:58]
  wire  a_sel_236 = _a_sel_T[236]; // @[ToAXI4.scala 242:58]
  wire  a_sel_237 = _a_sel_T[237]; // @[ToAXI4.scala 242:58]
  wire  a_sel_238 = _a_sel_T[238]; // @[ToAXI4.scala 242:58]
  wire  a_sel_239 = _a_sel_T[239]; // @[ToAXI4.scala 242:58]
  wire  a_sel_240 = _a_sel_T[240]; // @[ToAXI4.scala 242:58]
  wire  a_sel_241 = _a_sel_T[241]; // @[ToAXI4.scala 242:58]
  wire  a_sel_242 = _a_sel_T[242]; // @[ToAXI4.scala 242:58]
  wire  a_sel_243 = _a_sel_T[243]; // @[ToAXI4.scala 242:58]
  wire  a_sel_244 = _a_sel_T[244]; // @[ToAXI4.scala 242:58]
  wire  a_sel_245 = _a_sel_T[245]; // @[ToAXI4.scala 242:58]
  wire  a_sel_246 = _a_sel_T[246]; // @[ToAXI4.scala 242:58]
  wire  a_sel_247 = _a_sel_T[247]; // @[ToAXI4.scala 242:58]
  wire  a_sel_248 = _a_sel_T[248]; // @[ToAXI4.scala 242:58]
  wire  a_sel_249 = _a_sel_T[249]; // @[ToAXI4.scala 242:58]
  wire  a_sel_250 = _a_sel_T[250]; // @[ToAXI4.scala 242:58]
  wire  a_sel_251 = _a_sel_T[251]; // @[ToAXI4.scala 242:58]
  wire  a_sel_252 = _a_sel_T[252]; // @[ToAXI4.scala 242:58]
  wire  a_sel_253 = _a_sel_T[253]; // @[ToAXI4.scala 242:58]
  wire  a_sel_254 = _a_sel_T[254]; // @[ToAXI4.scala 242:58]
  wire  a_sel_255 = _a_sel_T[255]; // @[ToAXI4.scala 242:58]
  wire  a_sel_256 = _a_sel_T[256]; // @[ToAXI4.scala 242:58]
  wire  a_sel_257 = _a_sel_T[257]; // @[ToAXI4.scala 242:58]
  wire  a_sel_258 = _a_sel_T[258]; // @[ToAXI4.scala 242:58]
  wire  a_sel_259 = _a_sel_T[259]; // @[ToAXI4.scala 242:58]
  wire  a_sel_260 = _a_sel_T[260]; // @[ToAXI4.scala 242:58]
  wire  a_sel_261 = _a_sel_T[261]; // @[ToAXI4.scala 242:58]
  wire  a_sel_262 = _a_sel_T[262]; // @[ToAXI4.scala 242:58]
  wire  a_sel_263 = _a_sel_T[263]; // @[ToAXI4.scala 242:58]
  wire  a_sel_264 = _a_sel_T[264]; // @[ToAXI4.scala 242:58]
  wire  a_sel_265 = _a_sel_T[265]; // @[ToAXI4.scala 242:58]
  wire  a_sel_266 = _a_sel_T[266]; // @[ToAXI4.scala 242:58]
  wire  a_sel_267 = _a_sel_T[267]; // @[ToAXI4.scala 242:58]
  wire  a_sel_268 = _a_sel_T[268]; // @[ToAXI4.scala 242:58]
  wire  a_sel_269 = _a_sel_T[269]; // @[ToAXI4.scala 242:58]
  wire  a_sel_270 = _a_sel_T[270]; // @[ToAXI4.scala 242:58]
  wire  a_sel_271 = _a_sel_T[271]; // @[ToAXI4.scala 242:58]
  wire  a_sel_272 = _a_sel_T[272]; // @[ToAXI4.scala 242:58]
  wire  a_sel_273 = _a_sel_T[273]; // @[ToAXI4.scala 242:58]
  wire  a_sel_274 = _a_sel_T[274]; // @[ToAXI4.scala 242:58]
  wire  a_sel_275 = _a_sel_T[275]; // @[ToAXI4.scala 242:58]
  wire  a_sel_276 = _a_sel_T[276]; // @[ToAXI4.scala 242:58]
  wire  a_sel_277 = _a_sel_T[277]; // @[ToAXI4.scala 242:58]
  wire  a_sel_278 = _a_sel_T[278]; // @[ToAXI4.scala 242:58]
  wire  a_sel_279 = _a_sel_T[279]; // @[ToAXI4.scala 242:58]
  wire  a_sel_280 = _a_sel_T[280]; // @[ToAXI4.scala 242:58]
  wire  a_sel_281 = _a_sel_T[281]; // @[ToAXI4.scala 242:58]
  wire  a_sel_282 = _a_sel_T[282]; // @[ToAXI4.scala 242:58]
  wire  a_sel_283 = _a_sel_T[283]; // @[ToAXI4.scala 242:58]
  wire  a_sel_284 = _a_sel_T[284]; // @[ToAXI4.scala 242:58]
  wire  a_sel_285 = _a_sel_T[285]; // @[ToAXI4.scala 242:58]
  wire  a_sel_286 = _a_sel_T[286]; // @[ToAXI4.scala 242:58]
  wire  a_sel_287 = _a_sel_T[287]; // @[ToAXI4.scala 242:58]
  wire  a_sel_288 = _a_sel_T[288]; // @[ToAXI4.scala 242:58]
  wire  a_sel_289 = _a_sel_T[289]; // @[ToAXI4.scala 242:58]
  wire  a_sel_290 = _a_sel_T[290]; // @[ToAXI4.scala 242:58]
  wire  a_sel_291 = _a_sel_T[291]; // @[ToAXI4.scala 242:58]
  wire  a_sel_292 = _a_sel_T[292]; // @[ToAXI4.scala 242:58]
  wire  a_sel_293 = _a_sel_T[293]; // @[ToAXI4.scala 242:58]
  wire  a_sel_294 = _a_sel_T[294]; // @[ToAXI4.scala 242:58]
  wire  a_sel_295 = _a_sel_T[295]; // @[ToAXI4.scala 242:58]
  wire  a_sel_296 = _a_sel_T[296]; // @[ToAXI4.scala 242:58]
  wire  a_sel_297 = _a_sel_T[297]; // @[ToAXI4.scala 242:58]
  wire  a_sel_298 = _a_sel_T[298]; // @[ToAXI4.scala 242:58]
  wire  a_sel_299 = _a_sel_T[299]; // @[ToAXI4.scala 242:58]
  wire  a_sel_300 = _a_sel_T[300]; // @[ToAXI4.scala 242:58]
  wire  a_sel_301 = _a_sel_T[301]; // @[ToAXI4.scala 242:58]
  wire  a_sel_302 = _a_sel_T[302]; // @[ToAXI4.scala 242:58]
  wire  a_sel_303 = _a_sel_T[303]; // @[ToAXI4.scala 242:58]
  wire  a_sel_304 = _a_sel_T[304]; // @[ToAXI4.scala 242:58]
  wire  a_sel_305 = _a_sel_T[305]; // @[ToAXI4.scala 242:58]
  wire  a_sel_306 = _a_sel_T[306]; // @[ToAXI4.scala 242:58]
  wire  a_sel_307 = _a_sel_T[307]; // @[ToAXI4.scala 242:58]
  wire  a_sel_308 = _a_sel_T[308]; // @[ToAXI4.scala 242:58]
  wire  a_sel_309 = _a_sel_T[309]; // @[ToAXI4.scala 242:58]
  wire  a_sel_310 = _a_sel_T[310]; // @[ToAXI4.scala 242:58]
  wire  a_sel_311 = _a_sel_T[311]; // @[ToAXI4.scala 242:58]
  wire  a_sel_312 = _a_sel_T[312]; // @[ToAXI4.scala 242:58]
  wire  a_sel_313 = _a_sel_T[313]; // @[ToAXI4.scala 242:58]
  wire  a_sel_314 = _a_sel_T[314]; // @[ToAXI4.scala 242:58]
  wire  a_sel_315 = _a_sel_T[315]; // @[ToAXI4.scala 242:58]
  wire  a_sel_316 = _a_sel_T[316]; // @[ToAXI4.scala 242:58]
  wire  a_sel_317 = _a_sel_T[317]; // @[ToAXI4.scala 242:58]
  wire  a_sel_318 = _a_sel_T[318]; // @[ToAXI4.scala 242:58]
  wire  a_sel_319 = _a_sel_T[319]; // @[ToAXI4.scala 242:58]
  wire  a_sel_320 = _a_sel_T[320]; // @[ToAXI4.scala 242:58]
  wire  a_sel_321 = _a_sel_T[321]; // @[ToAXI4.scala 242:58]
  wire  a_sel_322 = _a_sel_T[322]; // @[ToAXI4.scala 242:58]
  wire  a_sel_323 = _a_sel_T[323]; // @[ToAXI4.scala 242:58]
  wire  a_sel_324 = _a_sel_T[324]; // @[ToAXI4.scala 242:58]
  wire  a_sel_325 = _a_sel_T[325]; // @[ToAXI4.scala 242:58]
  wire  a_sel_326 = _a_sel_T[326]; // @[ToAXI4.scala 242:58]
  wire  a_sel_327 = _a_sel_T[327]; // @[ToAXI4.scala 242:58]
  wire  a_sel_328 = _a_sel_T[328]; // @[ToAXI4.scala 242:58]
  wire  a_sel_329 = _a_sel_T[329]; // @[ToAXI4.scala 242:58]
  wire  a_sel_330 = _a_sel_T[330]; // @[ToAXI4.scala 242:58]
  wire  a_sel_331 = _a_sel_T[331]; // @[ToAXI4.scala 242:58]
  wire  a_sel_332 = _a_sel_T[332]; // @[ToAXI4.scala 242:58]
  wire  a_sel_333 = _a_sel_T[333]; // @[ToAXI4.scala 242:58]
  wire  a_sel_334 = _a_sel_T[334]; // @[ToAXI4.scala 242:58]
  wire  a_sel_335 = _a_sel_T[335]; // @[ToAXI4.scala 242:58]
  wire  a_sel_336 = _a_sel_T[336]; // @[ToAXI4.scala 242:58]
  wire  a_sel_337 = _a_sel_T[337]; // @[ToAXI4.scala 242:58]
  wire  a_sel_338 = _a_sel_T[338]; // @[ToAXI4.scala 242:58]
  wire  a_sel_339 = _a_sel_T[339]; // @[ToAXI4.scala 242:58]
  wire  a_sel_340 = _a_sel_T[340]; // @[ToAXI4.scala 242:58]
  wire  a_sel_341 = _a_sel_T[341]; // @[ToAXI4.scala 242:58]
  wire  a_sel_342 = _a_sel_T[342]; // @[ToAXI4.scala 242:58]
  wire  a_sel_343 = _a_sel_T[343]; // @[ToAXI4.scala 242:58]
  wire  a_sel_344 = _a_sel_T[344]; // @[ToAXI4.scala 242:58]
  wire  a_sel_345 = _a_sel_T[345]; // @[ToAXI4.scala 242:58]
  wire  a_sel_346 = _a_sel_T[346]; // @[ToAXI4.scala 242:58]
  wire  a_sel_347 = _a_sel_T[347]; // @[ToAXI4.scala 242:58]
  wire  a_sel_348 = _a_sel_T[348]; // @[ToAXI4.scala 242:58]
  wire  a_sel_349 = _a_sel_T[349]; // @[ToAXI4.scala 242:58]
  wire  a_sel_350 = _a_sel_T[350]; // @[ToAXI4.scala 242:58]
  wire  a_sel_351 = _a_sel_T[351]; // @[ToAXI4.scala 242:58]
  wire  a_sel_352 = _a_sel_T[352]; // @[ToAXI4.scala 242:58]
  wire  a_sel_353 = _a_sel_T[353]; // @[ToAXI4.scala 242:58]
  wire  a_sel_354 = _a_sel_T[354]; // @[ToAXI4.scala 242:58]
  wire  a_sel_355 = _a_sel_T[355]; // @[ToAXI4.scala 242:58]
  wire  a_sel_356 = _a_sel_T[356]; // @[ToAXI4.scala 242:58]
  wire  a_sel_357 = _a_sel_T[357]; // @[ToAXI4.scala 242:58]
  wire  a_sel_358 = _a_sel_T[358]; // @[ToAXI4.scala 242:58]
  wire  a_sel_359 = _a_sel_T[359]; // @[ToAXI4.scala 242:58]
  wire  a_sel_360 = _a_sel_T[360]; // @[ToAXI4.scala 242:58]
  wire  a_sel_361 = _a_sel_T[361]; // @[ToAXI4.scala 242:58]
  wire  a_sel_362 = _a_sel_T[362]; // @[ToAXI4.scala 242:58]
  wire  a_sel_363 = _a_sel_T[363]; // @[ToAXI4.scala 242:58]
  wire  a_sel_364 = _a_sel_T[364]; // @[ToAXI4.scala 242:58]
  wire  a_sel_365 = _a_sel_T[365]; // @[ToAXI4.scala 242:58]
  wire  a_sel_366 = _a_sel_T[366]; // @[ToAXI4.scala 242:58]
  wire  a_sel_367 = _a_sel_T[367]; // @[ToAXI4.scala 242:58]
  wire  a_sel_368 = _a_sel_T[368]; // @[ToAXI4.scala 242:58]
  wire  a_sel_369 = _a_sel_T[369]; // @[ToAXI4.scala 242:58]
  wire  a_sel_370 = _a_sel_T[370]; // @[ToAXI4.scala 242:58]
  wire  a_sel_371 = _a_sel_T[371]; // @[ToAXI4.scala 242:58]
  wire  a_sel_372 = _a_sel_T[372]; // @[ToAXI4.scala 242:58]
  wire  a_sel_373 = _a_sel_T[373]; // @[ToAXI4.scala 242:58]
  wire  a_sel_374 = _a_sel_T[374]; // @[ToAXI4.scala 242:58]
  wire  a_sel_375 = _a_sel_T[375]; // @[ToAXI4.scala 242:58]
  wire  a_sel_376 = _a_sel_T[376]; // @[ToAXI4.scala 242:58]
  wire  a_sel_377 = _a_sel_T[377]; // @[ToAXI4.scala 242:58]
  wire  a_sel_378 = _a_sel_T[378]; // @[ToAXI4.scala 242:58]
  wire  a_sel_379 = _a_sel_T[379]; // @[ToAXI4.scala 242:58]
  wire  a_sel_380 = _a_sel_T[380]; // @[ToAXI4.scala 242:58]
  wire  a_sel_381 = _a_sel_T[381]; // @[ToAXI4.scala 242:58]
  wire  a_sel_382 = _a_sel_T[382]; // @[ToAXI4.scala 242:58]
  wire  a_sel_383 = _a_sel_T[383]; // @[ToAXI4.scala 242:58]
  wire  a_sel_384 = _a_sel_T[384]; // @[ToAXI4.scala 242:58]
  wire  a_sel_385 = _a_sel_T[385]; // @[ToAXI4.scala 242:58]
  wire  a_sel_386 = _a_sel_T[386]; // @[ToAXI4.scala 242:58]
  wire  a_sel_387 = _a_sel_T[387]; // @[ToAXI4.scala 242:58]
  wire  a_sel_388 = _a_sel_T[388]; // @[ToAXI4.scala 242:58]
  wire  a_sel_389 = _a_sel_T[389]; // @[ToAXI4.scala 242:58]
  wire  a_sel_390 = _a_sel_T[390]; // @[ToAXI4.scala 242:58]
  wire  a_sel_391 = _a_sel_T[391]; // @[ToAXI4.scala 242:58]
  wire  a_sel_392 = _a_sel_T[392]; // @[ToAXI4.scala 242:58]
  wire  a_sel_393 = _a_sel_T[393]; // @[ToAXI4.scala 242:58]
  wire  a_sel_394 = _a_sel_T[394]; // @[ToAXI4.scala 242:58]
  wire  a_sel_395 = _a_sel_T[395]; // @[ToAXI4.scala 242:58]
  wire  a_sel_396 = _a_sel_T[396]; // @[ToAXI4.scala 242:58]
  wire  a_sel_397 = _a_sel_T[397]; // @[ToAXI4.scala 242:58]
  wire  a_sel_398 = _a_sel_T[398]; // @[ToAXI4.scala 242:58]
  wire  a_sel_399 = _a_sel_T[399]; // @[ToAXI4.scala 242:58]
  wire  a_sel_400 = _a_sel_T[400]; // @[ToAXI4.scala 242:58]
  wire  a_sel_401 = _a_sel_T[401]; // @[ToAXI4.scala 242:58]
  wire  a_sel_402 = _a_sel_T[402]; // @[ToAXI4.scala 242:58]
  wire  a_sel_403 = _a_sel_T[403]; // @[ToAXI4.scala 242:58]
  wire  a_sel_404 = _a_sel_T[404]; // @[ToAXI4.scala 242:58]
  wire  a_sel_405 = _a_sel_T[405]; // @[ToAXI4.scala 242:58]
  wire  a_sel_406 = _a_sel_T[406]; // @[ToAXI4.scala 242:58]
  wire  a_sel_407 = _a_sel_T[407]; // @[ToAXI4.scala 242:58]
  wire  a_sel_408 = _a_sel_T[408]; // @[ToAXI4.scala 242:58]
  wire  a_sel_409 = _a_sel_T[409]; // @[ToAXI4.scala 242:58]
  wire  a_sel_410 = _a_sel_T[410]; // @[ToAXI4.scala 242:58]
  wire  a_sel_411 = _a_sel_T[411]; // @[ToAXI4.scala 242:58]
  wire  a_sel_412 = _a_sel_T[412]; // @[ToAXI4.scala 242:58]
  wire  a_sel_413 = _a_sel_T[413]; // @[ToAXI4.scala 242:58]
  wire  a_sel_414 = _a_sel_T[414]; // @[ToAXI4.scala 242:58]
  wire  a_sel_415 = _a_sel_T[415]; // @[ToAXI4.scala 242:58]
  wire  a_sel_416 = _a_sel_T[416]; // @[ToAXI4.scala 242:58]
  wire  a_sel_417 = _a_sel_T[417]; // @[ToAXI4.scala 242:58]
  wire  a_sel_418 = _a_sel_T[418]; // @[ToAXI4.scala 242:58]
  wire  a_sel_419 = _a_sel_T[419]; // @[ToAXI4.scala 242:58]
  wire  a_sel_420 = _a_sel_T[420]; // @[ToAXI4.scala 242:58]
  wire  a_sel_421 = _a_sel_T[421]; // @[ToAXI4.scala 242:58]
  wire  a_sel_422 = _a_sel_T[422]; // @[ToAXI4.scala 242:58]
  wire  a_sel_423 = _a_sel_T[423]; // @[ToAXI4.scala 242:58]
  wire  a_sel_424 = _a_sel_T[424]; // @[ToAXI4.scala 242:58]
  wire  a_sel_425 = _a_sel_T[425]; // @[ToAXI4.scala 242:58]
  wire  a_sel_426 = _a_sel_T[426]; // @[ToAXI4.scala 242:58]
  wire  a_sel_427 = _a_sel_T[427]; // @[ToAXI4.scala 242:58]
  wire  a_sel_428 = _a_sel_T[428]; // @[ToAXI4.scala 242:58]
  wire  a_sel_429 = _a_sel_T[429]; // @[ToAXI4.scala 242:58]
  wire  a_sel_430 = _a_sel_T[430]; // @[ToAXI4.scala 242:58]
  wire  a_sel_431 = _a_sel_T[431]; // @[ToAXI4.scala 242:58]
  wire  a_sel_432 = _a_sel_T[432]; // @[ToAXI4.scala 242:58]
  wire  a_sel_433 = _a_sel_T[433]; // @[ToAXI4.scala 242:58]
  wire  a_sel_434 = _a_sel_T[434]; // @[ToAXI4.scala 242:58]
  wire  a_sel_435 = _a_sel_T[435]; // @[ToAXI4.scala 242:58]
  wire  a_sel_436 = _a_sel_T[436]; // @[ToAXI4.scala 242:58]
  wire  a_sel_437 = _a_sel_T[437]; // @[ToAXI4.scala 242:58]
  wire  a_sel_438 = _a_sel_T[438]; // @[ToAXI4.scala 242:58]
  wire  a_sel_439 = _a_sel_T[439]; // @[ToAXI4.scala 242:58]
  wire  a_sel_440 = _a_sel_T[440]; // @[ToAXI4.scala 242:58]
  wire  a_sel_441 = _a_sel_T[441]; // @[ToAXI4.scala 242:58]
  wire  a_sel_442 = _a_sel_T[442]; // @[ToAXI4.scala 242:58]
  wire  a_sel_443 = _a_sel_T[443]; // @[ToAXI4.scala 242:58]
  wire  a_sel_444 = _a_sel_T[444]; // @[ToAXI4.scala 242:58]
  wire  a_sel_445 = _a_sel_T[445]; // @[ToAXI4.scala 242:58]
  wire  a_sel_446 = _a_sel_T[446]; // @[ToAXI4.scala 242:58]
  wire  a_sel_447 = _a_sel_T[447]; // @[ToAXI4.scala 242:58]
  wire  a_sel_448 = _a_sel_T[448]; // @[ToAXI4.scala 242:58]
  wire  a_sel_449 = _a_sel_T[449]; // @[ToAXI4.scala 242:58]
  wire  a_sel_450 = _a_sel_T[450]; // @[ToAXI4.scala 242:58]
  wire  a_sel_451 = _a_sel_T[451]; // @[ToAXI4.scala 242:58]
  wire  a_sel_452 = _a_sel_T[452]; // @[ToAXI4.scala 242:58]
  wire  a_sel_453 = _a_sel_T[453]; // @[ToAXI4.scala 242:58]
  wire  a_sel_454 = _a_sel_T[454]; // @[ToAXI4.scala 242:58]
  wire  a_sel_455 = _a_sel_T[455]; // @[ToAXI4.scala 242:58]
  wire  a_sel_456 = _a_sel_T[456]; // @[ToAXI4.scala 242:58]
  wire  a_sel_457 = _a_sel_T[457]; // @[ToAXI4.scala 242:58]
  wire  a_sel_458 = _a_sel_T[458]; // @[ToAXI4.scala 242:58]
  wire  a_sel_459 = _a_sel_T[459]; // @[ToAXI4.scala 242:58]
  wire  a_sel_460 = _a_sel_T[460]; // @[ToAXI4.scala 242:58]
  wire  a_sel_461 = _a_sel_T[461]; // @[ToAXI4.scala 242:58]
  wire  a_sel_462 = _a_sel_T[462]; // @[ToAXI4.scala 242:58]
  wire  a_sel_463 = _a_sel_T[463]; // @[ToAXI4.scala 242:58]
  wire  a_sel_464 = _a_sel_T[464]; // @[ToAXI4.scala 242:58]
  wire  a_sel_465 = _a_sel_T[465]; // @[ToAXI4.scala 242:58]
  wire  a_sel_466 = _a_sel_T[466]; // @[ToAXI4.scala 242:58]
  wire  a_sel_467 = _a_sel_T[467]; // @[ToAXI4.scala 242:58]
  wire  a_sel_468 = _a_sel_T[468]; // @[ToAXI4.scala 242:58]
  wire  a_sel_469 = _a_sel_T[469]; // @[ToAXI4.scala 242:58]
  wire  a_sel_470 = _a_sel_T[470]; // @[ToAXI4.scala 242:58]
  wire  a_sel_471 = _a_sel_T[471]; // @[ToAXI4.scala 242:58]
  wire  a_sel_472 = _a_sel_T[472]; // @[ToAXI4.scala 242:58]
  wire  a_sel_473 = _a_sel_T[473]; // @[ToAXI4.scala 242:58]
  wire  a_sel_474 = _a_sel_T[474]; // @[ToAXI4.scala 242:58]
  wire  a_sel_475 = _a_sel_T[475]; // @[ToAXI4.scala 242:58]
  wire  a_sel_476 = _a_sel_T[476]; // @[ToAXI4.scala 242:58]
  wire  a_sel_477 = _a_sel_T[477]; // @[ToAXI4.scala 242:58]
  wire  a_sel_478 = _a_sel_T[478]; // @[ToAXI4.scala 242:58]
  wire  a_sel_479 = _a_sel_T[479]; // @[ToAXI4.scala 242:58]
  wire  a_sel_480 = _a_sel_T[480]; // @[ToAXI4.scala 242:58]
  wire  a_sel_481 = _a_sel_T[481]; // @[ToAXI4.scala 242:58]
  wire  a_sel_482 = _a_sel_T[482]; // @[ToAXI4.scala 242:58]
  wire  a_sel_483 = _a_sel_T[483]; // @[ToAXI4.scala 242:58]
  wire  a_sel_484 = _a_sel_T[484]; // @[ToAXI4.scala 242:58]
  wire  a_sel_485 = _a_sel_T[485]; // @[ToAXI4.scala 242:58]
  wire  a_sel_486 = _a_sel_T[486]; // @[ToAXI4.scala 242:58]
  wire  a_sel_487 = _a_sel_T[487]; // @[ToAXI4.scala 242:58]
  wire  a_sel_488 = _a_sel_T[488]; // @[ToAXI4.scala 242:58]
  wire  a_sel_489 = _a_sel_T[489]; // @[ToAXI4.scala 242:58]
  wire  a_sel_490 = _a_sel_T[490]; // @[ToAXI4.scala 242:58]
  wire  a_sel_491 = _a_sel_T[491]; // @[ToAXI4.scala 242:58]
  wire  a_sel_492 = _a_sel_T[492]; // @[ToAXI4.scala 242:58]
  wire  a_sel_493 = _a_sel_T[493]; // @[ToAXI4.scala 242:58]
  wire  a_sel_494 = _a_sel_T[494]; // @[ToAXI4.scala 242:58]
  wire  a_sel_495 = _a_sel_T[495]; // @[ToAXI4.scala 242:58]
  wire  a_sel_496 = _a_sel_T[496]; // @[ToAXI4.scala 242:58]
  wire  a_sel_497 = _a_sel_T[497]; // @[ToAXI4.scala 242:58]
  wire  a_sel_498 = _a_sel_T[498]; // @[ToAXI4.scala 242:58]
  wire  a_sel_499 = _a_sel_T[499]; // @[ToAXI4.scala 242:58]
  wire  a_sel_500 = _a_sel_T[500]; // @[ToAXI4.scala 242:58]
  wire  a_sel_501 = _a_sel_T[501]; // @[ToAXI4.scala 242:58]
  wire  a_sel_502 = _a_sel_T[502]; // @[ToAXI4.scala 242:58]
  wire  a_sel_503 = _a_sel_T[503]; // @[ToAXI4.scala 242:58]
  wire  a_sel_504 = _a_sel_T[504]; // @[ToAXI4.scala 242:58]
  wire  a_sel_505 = _a_sel_T[505]; // @[ToAXI4.scala 242:58]
  wire  a_sel_506 = _a_sel_T[506]; // @[ToAXI4.scala 242:58]
  wire  a_sel_507 = _a_sel_T[507]; // @[ToAXI4.scala 242:58]
  wire  a_sel_508 = _a_sel_T[508]; // @[ToAXI4.scala 242:58]
  wire  a_sel_509 = _a_sel_T[509]; // @[ToAXI4.scala 242:58]
  wire  a_sel_510 = _a_sel_T[510]; // @[ToAXI4.scala 242:58]
  wire  a_sel_511 = _a_sel_T[511]; // @[ToAXI4.scala 242:58]
  wire [8:0] d_sel_shiftAmount = r_wins ? auto_out_r_bits_id : auto_out_b_bits_id; // @[ToAXI4.scala 243:31]
  wire [511:0] _d_sel_T_1 = 512'h1 << d_sel_shiftAmount; // @[OneHot.scala 64:12]
  wire  d_sel_0 = _d_sel_T_1[0]; // @[ToAXI4.scala 243:93]
  wire  d_sel_1 = _d_sel_T_1[1]; // @[ToAXI4.scala 243:93]
  wire  d_sel_2 = _d_sel_T_1[2]; // @[ToAXI4.scala 243:93]
  wire  d_sel_3 = _d_sel_T_1[3]; // @[ToAXI4.scala 243:93]
  wire  d_sel_4 = _d_sel_T_1[4]; // @[ToAXI4.scala 243:93]
  wire  d_sel_5 = _d_sel_T_1[5]; // @[ToAXI4.scala 243:93]
  wire  d_sel_6 = _d_sel_T_1[6]; // @[ToAXI4.scala 243:93]
  wire  d_sel_7 = _d_sel_T_1[7]; // @[ToAXI4.scala 243:93]
  wire  d_sel_8 = _d_sel_T_1[8]; // @[ToAXI4.scala 243:93]
  wire  d_sel_9 = _d_sel_T_1[9]; // @[ToAXI4.scala 243:93]
  wire  d_sel_10 = _d_sel_T_1[10]; // @[ToAXI4.scala 243:93]
  wire  d_sel_11 = _d_sel_T_1[11]; // @[ToAXI4.scala 243:93]
  wire  d_sel_12 = _d_sel_T_1[12]; // @[ToAXI4.scala 243:93]
  wire  d_sel_13 = _d_sel_T_1[13]; // @[ToAXI4.scala 243:93]
  wire  d_sel_14 = _d_sel_T_1[14]; // @[ToAXI4.scala 243:93]
  wire  d_sel_15 = _d_sel_T_1[15]; // @[ToAXI4.scala 243:93]
  wire  d_sel_16 = _d_sel_T_1[16]; // @[ToAXI4.scala 243:93]
  wire  d_sel_17 = _d_sel_T_1[17]; // @[ToAXI4.scala 243:93]
  wire  d_sel_18 = _d_sel_T_1[18]; // @[ToAXI4.scala 243:93]
  wire  d_sel_19 = _d_sel_T_1[19]; // @[ToAXI4.scala 243:93]
  wire  d_sel_20 = _d_sel_T_1[20]; // @[ToAXI4.scala 243:93]
  wire  d_sel_21 = _d_sel_T_1[21]; // @[ToAXI4.scala 243:93]
  wire  d_sel_22 = _d_sel_T_1[22]; // @[ToAXI4.scala 243:93]
  wire  d_sel_23 = _d_sel_T_1[23]; // @[ToAXI4.scala 243:93]
  wire  d_sel_24 = _d_sel_T_1[24]; // @[ToAXI4.scala 243:93]
  wire  d_sel_25 = _d_sel_T_1[25]; // @[ToAXI4.scala 243:93]
  wire  d_sel_26 = _d_sel_T_1[26]; // @[ToAXI4.scala 243:93]
  wire  d_sel_27 = _d_sel_T_1[27]; // @[ToAXI4.scala 243:93]
  wire  d_sel_28 = _d_sel_T_1[28]; // @[ToAXI4.scala 243:93]
  wire  d_sel_29 = _d_sel_T_1[29]; // @[ToAXI4.scala 243:93]
  wire  d_sel_30 = _d_sel_T_1[30]; // @[ToAXI4.scala 243:93]
  wire  d_sel_31 = _d_sel_T_1[31]; // @[ToAXI4.scala 243:93]
  wire  d_sel_32 = _d_sel_T_1[32]; // @[ToAXI4.scala 243:93]
  wire  d_sel_33 = _d_sel_T_1[33]; // @[ToAXI4.scala 243:93]
  wire  d_sel_34 = _d_sel_T_1[34]; // @[ToAXI4.scala 243:93]
  wire  d_sel_35 = _d_sel_T_1[35]; // @[ToAXI4.scala 243:93]
  wire  d_sel_36 = _d_sel_T_1[36]; // @[ToAXI4.scala 243:93]
  wire  d_sel_37 = _d_sel_T_1[37]; // @[ToAXI4.scala 243:93]
  wire  d_sel_38 = _d_sel_T_1[38]; // @[ToAXI4.scala 243:93]
  wire  d_sel_39 = _d_sel_T_1[39]; // @[ToAXI4.scala 243:93]
  wire  d_sel_40 = _d_sel_T_1[40]; // @[ToAXI4.scala 243:93]
  wire  d_sel_41 = _d_sel_T_1[41]; // @[ToAXI4.scala 243:93]
  wire  d_sel_42 = _d_sel_T_1[42]; // @[ToAXI4.scala 243:93]
  wire  d_sel_43 = _d_sel_T_1[43]; // @[ToAXI4.scala 243:93]
  wire  d_sel_44 = _d_sel_T_1[44]; // @[ToAXI4.scala 243:93]
  wire  d_sel_45 = _d_sel_T_1[45]; // @[ToAXI4.scala 243:93]
  wire  d_sel_46 = _d_sel_T_1[46]; // @[ToAXI4.scala 243:93]
  wire  d_sel_47 = _d_sel_T_1[47]; // @[ToAXI4.scala 243:93]
  wire  d_sel_48 = _d_sel_T_1[48]; // @[ToAXI4.scala 243:93]
  wire  d_sel_49 = _d_sel_T_1[49]; // @[ToAXI4.scala 243:93]
  wire  d_sel_50 = _d_sel_T_1[50]; // @[ToAXI4.scala 243:93]
  wire  d_sel_51 = _d_sel_T_1[51]; // @[ToAXI4.scala 243:93]
  wire  d_sel_52 = _d_sel_T_1[52]; // @[ToAXI4.scala 243:93]
  wire  d_sel_53 = _d_sel_T_1[53]; // @[ToAXI4.scala 243:93]
  wire  d_sel_54 = _d_sel_T_1[54]; // @[ToAXI4.scala 243:93]
  wire  d_sel_55 = _d_sel_T_1[55]; // @[ToAXI4.scala 243:93]
  wire  d_sel_56 = _d_sel_T_1[56]; // @[ToAXI4.scala 243:93]
  wire  d_sel_57 = _d_sel_T_1[57]; // @[ToAXI4.scala 243:93]
  wire  d_sel_58 = _d_sel_T_1[58]; // @[ToAXI4.scala 243:93]
  wire  d_sel_59 = _d_sel_T_1[59]; // @[ToAXI4.scala 243:93]
  wire  d_sel_60 = _d_sel_T_1[60]; // @[ToAXI4.scala 243:93]
  wire  d_sel_61 = _d_sel_T_1[61]; // @[ToAXI4.scala 243:93]
  wire  d_sel_62 = _d_sel_T_1[62]; // @[ToAXI4.scala 243:93]
  wire  d_sel_63 = _d_sel_T_1[63]; // @[ToAXI4.scala 243:93]
  wire  d_sel_64 = _d_sel_T_1[64]; // @[ToAXI4.scala 243:93]
  wire  d_sel_65 = _d_sel_T_1[65]; // @[ToAXI4.scala 243:93]
  wire  d_sel_66 = _d_sel_T_1[66]; // @[ToAXI4.scala 243:93]
  wire  d_sel_67 = _d_sel_T_1[67]; // @[ToAXI4.scala 243:93]
  wire  d_sel_68 = _d_sel_T_1[68]; // @[ToAXI4.scala 243:93]
  wire  d_sel_69 = _d_sel_T_1[69]; // @[ToAXI4.scala 243:93]
  wire  d_sel_70 = _d_sel_T_1[70]; // @[ToAXI4.scala 243:93]
  wire  d_sel_71 = _d_sel_T_1[71]; // @[ToAXI4.scala 243:93]
  wire  d_sel_72 = _d_sel_T_1[72]; // @[ToAXI4.scala 243:93]
  wire  d_sel_73 = _d_sel_T_1[73]; // @[ToAXI4.scala 243:93]
  wire  d_sel_74 = _d_sel_T_1[74]; // @[ToAXI4.scala 243:93]
  wire  d_sel_75 = _d_sel_T_1[75]; // @[ToAXI4.scala 243:93]
  wire  d_sel_76 = _d_sel_T_1[76]; // @[ToAXI4.scala 243:93]
  wire  d_sel_77 = _d_sel_T_1[77]; // @[ToAXI4.scala 243:93]
  wire  d_sel_78 = _d_sel_T_1[78]; // @[ToAXI4.scala 243:93]
  wire  d_sel_79 = _d_sel_T_1[79]; // @[ToAXI4.scala 243:93]
  wire  d_sel_80 = _d_sel_T_1[80]; // @[ToAXI4.scala 243:93]
  wire  d_sel_81 = _d_sel_T_1[81]; // @[ToAXI4.scala 243:93]
  wire  d_sel_82 = _d_sel_T_1[82]; // @[ToAXI4.scala 243:93]
  wire  d_sel_83 = _d_sel_T_1[83]; // @[ToAXI4.scala 243:93]
  wire  d_sel_84 = _d_sel_T_1[84]; // @[ToAXI4.scala 243:93]
  wire  d_sel_85 = _d_sel_T_1[85]; // @[ToAXI4.scala 243:93]
  wire  d_sel_86 = _d_sel_T_1[86]; // @[ToAXI4.scala 243:93]
  wire  d_sel_87 = _d_sel_T_1[87]; // @[ToAXI4.scala 243:93]
  wire  d_sel_88 = _d_sel_T_1[88]; // @[ToAXI4.scala 243:93]
  wire  d_sel_89 = _d_sel_T_1[89]; // @[ToAXI4.scala 243:93]
  wire  d_sel_90 = _d_sel_T_1[90]; // @[ToAXI4.scala 243:93]
  wire  d_sel_91 = _d_sel_T_1[91]; // @[ToAXI4.scala 243:93]
  wire  d_sel_92 = _d_sel_T_1[92]; // @[ToAXI4.scala 243:93]
  wire  d_sel_93 = _d_sel_T_1[93]; // @[ToAXI4.scala 243:93]
  wire  d_sel_94 = _d_sel_T_1[94]; // @[ToAXI4.scala 243:93]
  wire  d_sel_95 = _d_sel_T_1[95]; // @[ToAXI4.scala 243:93]
  wire  d_sel_96 = _d_sel_T_1[96]; // @[ToAXI4.scala 243:93]
  wire  d_sel_97 = _d_sel_T_1[97]; // @[ToAXI4.scala 243:93]
  wire  d_sel_98 = _d_sel_T_1[98]; // @[ToAXI4.scala 243:93]
  wire  d_sel_99 = _d_sel_T_1[99]; // @[ToAXI4.scala 243:93]
  wire  d_sel_100 = _d_sel_T_1[100]; // @[ToAXI4.scala 243:93]
  wire  d_sel_101 = _d_sel_T_1[101]; // @[ToAXI4.scala 243:93]
  wire  d_sel_102 = _d_sel_T_1[102]; // @[ToAXI4.scala 243:93]
  wire  d_sel_103 = _d_sel_T_1[103]; // @[ToAXI4.scala 243:93]
  wire  d_sel_104 = _d_sel_T_1[104]; // @[ToAXI4.scala 243:93]
  wire  d_sel_105 = _d_sel_T_1[105]; // @[ToAXI4.scala 243:93]
  wire  d_sel_106 = _d_sel_T_1[106]; // @[ToAXI4.scala 243:93]
  wire  d_sel_107 = _d_sel_T_1[107]; // @[ToAXI4.scala 243:93]
  wire  d_sel_108 = _d_sel_T_1[108]; // @[ToAXI4.scala 243:93]
  wire  d_sel_109 = _d_sel_T_1[109]; // @[ToAXI4.scala 243:93]
  wire  d_sel_110 = _d_sel_T_1[110]; // @[ToAXI4.scala 243:93]
  wire  d_sel_111 = _d_sel_T_1[111]; // @[ToAXI4.scala 243:93]
  wire  d_sel_112 = _d_sel_T_1[112]; // @[ToAXI4.scala 243:93]
  wire  d_sel_113 = _d_sel_T_1[113]; // @[ToAXI4.scala 243:93]
  wire  d_sel_114 = _d_sel_T_1[114]; // @[ToAXI4.scala 243:93]
  wire  d_sel_115 = _d_sel_T_1[115]; // @[ToAXI4.scala 243:93]
  wire  d_sel_116 = _d_sel_T_1[116]; // @[ToAXI4.scala 243:93]
  wire  d_sel_117 = _d_sel_T_1[117]; // @[ToAXI4.scala 243:93]
  wire  d_sel_118 = _d_sel_T_1[118]; // @[ToAXI4.scala 243:93]
  wire  d_sel_119 = _d_sel_T_1[119]; // @[ToAXI4.scala 243:93]
  wire  d_sel_120 = _d_sel_T_1[120]; // @[ToAXI4.scala 243:93]
  wire  d_sel_121 = _d_sel_T_1[121]; // @[ToAXI4.scala 243:93]
  wire  d_sel_122 = _d_sel_T_1[122]; // @[ToAXI4.scala 243:93]
  wire  d_sel_123 = _d_sel_T_1[123]; // @[ToAXI4.scala 243:93]
  wire  d_sel_124 = _d_sel_T_1[124]; // @[ToAXI4.scala 243:93]
  wire  d_sel_125 = _d_sel_T_1[125]; // @[ToAXI4.scala 243:93]
  wire  d_sel_126 = _d_sel_T_1[126]; // @[ToAXI4.scala 243:93]
  wire  d_sel_127 = _d_sel_T_1[127]; // @[ToAXI4.scala 243:93]
  wire  d_sel_128 = _d_sel_T_1[128]; // @[ToAXI4.scala 243:93]
  wire  d_sel_129 = _d_sel_T_1[129]; // @[ToAXI4.scala 243:93]
  wire  d_sel_130 = _d_sel_T_1[130]; // @[ToAXI4.scala 243:93]
  wire  d_sel_131 = _d_sel_T_1[131]; // @[ToAXI4.scala 243:93]
  wire  d_sel_132 = _d_sel_T_1[132]; // @[ToAXI4.scala 243:93]
  wire  d_sel_133 = _d_sel_T_1[133]; // @[ToAXI4.scala 243:93]
  wire  d_sel_134 = _d_sel_T_1[134]; // @[ToAXI4.scala 243:93]
  wire  d_sel_135 = _d_sel_T_1[135]; // @[ToAXI4.scala 243:93]
  wire  d_sel_136 = _d_sel_T_1[136]; // @[ToAXI4.scala 243:93]
  wire  d_sel_137 = _d_sel_T_1[137]; // @[ToAXI4.scala 243:93]
  wire  d_sel_138 = _d_sel_T_1[138]; // @[ToAXI4.scala 243:93]
  wire  d_sel_139 = _d_sel_T_1[139]; // @[ToAXI4.scala 243:93]
  wire  d_sel_140 = _d_sel_T_1[140]; // @[ToAXI4.scala 243:93]
  wire  d_sel_141 = _d_sel_T_1[141]; // @[ToAXI4.scala 243:93]
  wire  d_sel_142 = _d_sel_T_1[142]; // @[ToAXI4.scala 243:93]
  wire  d_sel_143 = _d_sel_T_1[143]; // @[ToAXI4.scala 243:93]
  wire  d_sel_144 = _d_sel_T_1[144]; // @[ToAXI4.scala 243:93]
  wire  d_sel_145 = _d_sel_T_1[145]; // @[ToAXI4.scala 243:93]
  wire  d_sel_146 = _d_sel_T_1[146]; // @[ToAXI4.scala 243:93]
  wire  d_sel_147 = _d_sel_T_1[147]; // @[ToAXI4.scala 243:93]
  wire  d_sel_148 = _d_sel_T_1[148]; // @[ToAXI4.scala 243:93]
  wire  d_sel_149 = _d_sel_T_1[149]; // @[ToAXI4.scala 243:93]
  wire  d_sel_150 = _d_sel_T_1[150]; // @[ToAXI4.scala 243:93]
  wire  d_sel_151 = _d_sel_T_1[151]; // @[ToAXI4.scala 243:93]
  wire  d_sel_152 = _d_sel_T_1[152]; // @[ToAXI4.scala 243:93]
  wire  d_sel_153 = _d_sel_T_1[153]; // @[ToAXI4.scala 243:93]
  wire  d_sel_154 = _d_sel_T_1[154]; // @[ToAXI4.scala 243:93]
  wire  d_sel_155 = _d_sel_T_1[155]; // @[ToAXI4.scala 243:93]
  wire  d_sel_156 = _d_sel_T_1[156]; // @[ToAXI4.scala 243:93]
  wire  d_sel_157 = _d_sel_T_1[157]; // @[ToAXI4.scala 243:93]
  wire  d_sel_158 = _d_sel_T_1[158]; // @[ToAXI4.scala 243:93]
  wire  d_sel_159 = _d_sel_T_1[159]; // @[ToAXI4.scala 243:93]
  wire  d_sel_160 = _d_sel_T_1[160]; // @[ToAXI4.scala 243:93]
  wire  d_sel_161 = _d_sel_T_1[161]; // @[ToAXI4.scala 243:93]
  wire  d_sel_162 = _d_sel_T_1[162]; // @[ToAXI4.scala 243:93]
  wire  d_sel_163 = _d_sel_T_1[163]; // @[ToAXI4.scala 243:93]
  wire  d_sel_164 = _d_sel_T_1[164]; // @[ToAXI4.scala 243:93]
  wire  d_sel_165 = _d_sel_T_1[165]; // @[ToAXI4.scala 243:93]
  wire  d_sel_166 = _d_sel_T_1[166]; // @[ToAXI4.scala 243:93]
  wire  d_sel_167 = _d_sel_T_1[167]; // @[ToAXI4.scala 243:93]
  wire  d_sel_168 = _d_sel_T_1[168]; // @[ToAXI4.scala 243:93]
  wire  d_sel_169 = _d_sel_T_1[169]; // @[ToAXI4.scala 243:93]
  wire  d_sel_170 = _d_sel_T_1[170]; // @[ToAXI4.scala 243:93]
  wire  d_sel_171 = _d_sel_T_1[171]; // @[ToAXI4.scala 243:93]
  wire  d_sel_172 = _d_sel_T_1[172]; // @[ToAXI4.scala 243:93]
  wire  d_sel_173 = _d_sel_T_1[173]; // @[ToAXI4.scala 243:93]
  wire  d_sel_174 = _d_sel_T_1[174]; // @[ToAXI4.scala 243:93]
  wire  d_sel_175 = _d_sel_T_1[175]; // @[ToAXI4.scala 243:93]
  wire  d_sel_176 = _d_sel_T_1[176]; // @[ToAXI4.scala 243:93]
  wire  d_sel_177 = _d_sel_T_1[177]; // @[ToAXI4.scala 243:93]
  wire  d_sel_178 = _d_sel_T_1[178]; // @[ToAXI4.scala 243:93]
  wire  d_sel_179 = _d_sel_T_1[179]; // @[ToAXI4.scala 243:93]
  wire  d_sel_180 = _d_sel_T_1[180]; // @[ToAXI4.scala 243:93]
  wire  d_sel_181 = _d_sel_T_1[181]; // @[ToAXI4.scala 243:93]
  wire  d_sel_182 = _d_sel_T_1[182]; // @[ToAXI4.scala 243:93]
  wire  d_sel_183 = _d_sel_T_1[183]; // @[ToAXI4.scala 243:93]
  wire  d_sel_184 = _d_sel_T_1[184]; // @[ToAXI4.scala 243:93]
  wire  d_sel_185 = _d_sel_T_1[185]; // @[ToAXI4.scala 243:93]
  wire  d_sel_186 = _d_sel_T_1[186]; // @[ToAXI4.scala 243:93]
  wire  d_sel_187 = _d_sel_T_1[187]; // @[ToAXI4.scala 243:93]
  wire  d_sel_188 = _d_sel_T_1[188]; // @[ToAXI4.scala 243:93]
  wire  d_sel_189 = _d_sel_T_1[189]; // @[ToAXI4.scala 243:93]
  wire  d_sel_190 = _d_sel_T_1[190]; // @[ToAXI4.scala 243:93]
  wire  d_sel_191 = _d_sel_T_1[191]; // @[ToAXI4.scala 243:93]
  wire  d_sel_192 = _d_sel_T_1[192]; // @[ToAXI4.scala 243:93]
  wire  d_sel_193 = _d_sel_T_1[193]; // @[ToAXI4.scala 243:93]
  wire  d_sel_194 = _d_sel_T_1[194]; // @[ToAXI4.scala 243:93]
  wire  d_sel_195 = _d_sel_T_1[195]; // @[ToAXI4.scala 243:93]
  wire  d_sel_196 = _d_sel_T_1[196]; // @[ToAXI4.scala 243:93]
  wire  d_sel_197 = _d_sel_T_1[197]; // @[ToAXI4.scala 243:93]
  wire  d_sel_198 = _d_sel_T_1[198]; // @[ToAXI4.scala 243:93]
  wire  d_sel_199 = _d_sel_T_1[199]; // @[ToAXI4.scala 243:93]
  wire  d_sel_200 = _d_sel_T_1[200]; // @[ToAXI4.scala 243:93]
  wire  d_sel_201 = _d_sel_T_1[201]; // @[ToAXI4.scala 243:93]
  wire  d_sel_202 = _d_sel_T_1[202]; // @[ToAXI4.scala 243:93]
  wire  d_sel_203 = _d_sel_T_1[203]; // @[ToAXI4.scala 243:93]
  wire  d_sel_204 = _d_sel_T_1[204]; // @[ToAXI4.scala 243:93]
  wire  d_sel_205 = _d_sel_T_1[205]; // @[ToAXI4.scala 243:93]
  wire  d_sel_206 = _d_sel_T_1[206]; // @[ToAXI4.scala 243:93]
  wire  d_sel_207 = _d_sel_T_1[207]; // @[ToAXI4.scala 243:93]
  wire  d_sel_208 = _d_sel_T_1[208]; // @[ToAXI4.scala 243:93]
  wire  d_sel_209 = _d_sel_T_1[209]; // @[ToAXI4.scala 243:93]
  wire  d_sel_210 = _d_sel_T_1[210]; // @[ToAXI4.scala 243:93]
  wire  d_sel_211 = _d_sel_T_1[211]; // @[ToAXI4.scala 243:93]
  wire  d_sel_212 = _d_sel_T_1[212]; // @[ToAXI4.scala 243:93]
  wire  d_sel_213 = _d_sel_T_1[213]; // @[ToAXI4.scala 243:93]
  wire  d_sel_214 = _d_sel_T_1[214]; // @[ToAXI4.scala 243:93]
  wire  d_sel_215 = _d_sel_T_1[215]; // @[ToAXI4.scala 243:93]
  wire  d_sel_216 = _d_sel_T_1[216]; // @[ToAXI4.scala 243:93]
  wire  d_sel_217 = _d_sel_T_1[217]; // @[ToAXI4.scala 243:93]
  wire  d_sel_218 = _d_sel_T_1[218]; // @[ToAXI4.scala 243:93]
  wire  d_sel_219 = _d_sel_T_1[219]; // @[ToAXI4.scala 243:93]
  wire  d_sel_220 = _d_sel_T_1[220]; // @[ToAXI4.scala 243:93]
  wire  d_sel_221 = _d_sel_T_1[221]; // @[ToAXI4.scala 243:93]
  wire  d_sel_222 = _d_sel_T_1[222]; // @[ToAXI4.scala 243:93]
  wire  d_sel_223 = _d_sel_T_1[223]; // @[ToAXI4.scala 243:93]
  wire  d_sel_224 = _d_sel_T_1[224]; // @[ToAXI4.scala 243:93]
  wire  d_sel_225 = _d_sel_T_1[225]; // @[ToAXI4.scala 243:93]
  wire  d_sel_226 = _d_sel_T_1[226]; // @[ToAXI4.scala 243:93]
  wire  d_sel_227 = _d_sel_T_1[227]; // @[ToAXI4.scala 243:93]
  wire  d_sel_228 = _d_sel_T_1[228]; // @[ToAXI4.scala 243:93]
  wire  d_sel_229 = _d_sel_T_1[229]; // @[ToAXI4.scala 243:93]
  wire  d_sel_230 = _d_sel_T_1[230]; // @[ToAXI4.scala 243:93]
  wire  d_sel_231 = _d_sel_T_1[231]; // @[ToAXI4.scala 243:93]
  wire  d_sel_232 = _d_sel_T_1[232]; // @[ToAXI4.scala 243:93]
  wire  d_sel_233 = _d_sel_T_1[233]; // @[ToAXI4.scala 243:93]
  wire  d_sel_234 = _d_sel_T_1[234]; // @[ToAXI4.scala 243:93]
  wire  d_sel_235 = _d_sel_T_1[235]; // @[ToAXI4.scala 243:93]
  wire  d_sel_236 = _d_sel_T_1[236]; // @[ToAXI4.scala 243:93]
  wire  d_sel_237 = _d_sel_T_1[237]; // @[ToAXI4.scala 243:93]
  wire  d_sel_238 = _d_sel_T_1[238]; // @[ToAXI4.scala 243:93]
  wire  d_sel_239 = _d_sel_T_1[239]; // @[ToAXI4.scala 243:93]
  wire  d_sel_240 = _d_sel_T_1[240]; // @[ToAXI4.scala 243:93]
  wire  d_sel_241 = _d_sel_T_1[241]; // @[ToAXI4.scala 243:93]
  wire  d_sel_242 = _d_sel_T_1[242]; // @[ToAXI4.scala 243:93]
  wire  d_sel_243 = _d_sel_T_1[243]; // @[ToAXI4.scala 243:93]
  wire  d_sel_244 = _d_sel_T_1[244]; // @[ToAXI4.scala 243:93]
  wire  d_sel_245 = _d_sel_T_1[245]; // @[ToAXI4.scala 243:93]
  wire  d_sel_246 = _d_sel_T_1[246]; // @[ToAXI4.scala 243:93]
  wire  d_sel_247 = _d_sel_T_1[247]; // @[ToAXI4.scala 243:93]
  wire  d_sel_248 = _d_sel_T_1[248]; // @[ToAXI4.scala 243:93]
  wire  d_sel_249 = _d_sel_T_1[249]; // @[ToAXI4.scala 243:93]
  wire  d_sel_250 = _d_sel_T_1[250]; // @[ToAXI4.scala 243:93]
  wire  d_sel_251 = _d_sel_T_1[251]; // @[ToAXI4.scala 243:93]
  wire  d_sel_252 = _d_sel_T_1[252]; // @[ToAXI4.scala 243:93]
  wire  d_sel_253 = _d_sel_T_1[253]; // @[ToAXI4.scala 243:93]
  wire  d_sel_254 = _d_sel_T_1[254]; // @[ToAXI4.scala 243:93]
  wire  d_sel_255 = _d_sel_T_1[255]; // @[ToAXI4.scala 243:93]
  wire  d_sel_256 = _d_sel_T_1[256]; // @[ToAXI4.scala 243:93]
  wire  d_sel_257 = _d_sel_T_1[257]; // @[ToAXI4.scala 243:93]
  wire  d_sel_258 = _d_sel_T_1[258]; // @[ToAXI4.scala 243:93]
  wire  d_sel_259 = _d_sel_T_1[259]; // @[ToAXI4.scala 243:93]
  wire  d_sel_260 = _d_sel_T_1[260]; // @[ToAXI4.scala 243:93]
  wire  d_sel_261 = _d_sel_T_1[261]; // @[ToAXI4.scala 243:93]
  wire  d_sel_262 = _d_sel_T_1[262]; // @[ToAXI4.scala 243:93]
  wire  d_sel_263 = _d_sel_T_1[263]; // @[ToAXI4.scala 243:93]
  wire  d_sel_264 = _d_sel_T_1[264]; // @[ToAXI4.scala 243:93]
  wire  d_sel_265 = _d_sel_T_1[265]; // @[ToAXI4.scala 243:93]
  wire  d_sel_266 = _d_sel_T_1[266]; // @[ToAXI4.scala 243:93]
  wire  d_sel_267 = _d_sel_T_1[267]; // @[ToAXI4.scala 243:93]
  wire  d_sel_268 = _d_sel_T_1[268]; // @[ToAXI4.scala 243:93]
  wire  d_sel_269 = _d_sel_T_1[269]; // @[ToAXI4.scala 243:93]
  wire  d_sel_270 = _d_sel_T_1[270]; // @[ToAXI4.scala 243:93]
  wire  d_sel_271 = _d_sel_T_1[271]; // @[ToAXI4.scala 243:93]
  wire  d_sel_272 = _d_sel_T_1[272]; // @[ToAXI4.scala 243:93]
  wire  d_sel_273 = _d_sel_T_1[273]; // @[ToAXI4.scala 243:93]
  wire  d_sel_274 = _d_sel_T_1[274]; // @[ToAXI4.scala 243:93]
  wire  d_sel_275 = _d_sel_T_1[275]; // @[ToAXI4.scala 243:93]
  wire  d_sel_276 = _d_sel_T_1[276]; // @[ToAXI4.scala 243:93]
  wire  d_sel_277 = _d_sel_T_1[277]; // @[ToAXI4.scala 243:93]
  wire  d_sel_278 = _d_sel_T_1[278]; // @[ToAXI4.scala 243:93]
  wire  d_sel_279 = _d_sel_T_1[279]; // @[ToAXI4.scala 243:93]
  wire  d_sel_280 = _d_sel_T_1[280]; // @[ToAXI4.scala 243:93]
  wire  d_sel_281 = _d_sel_T_1[281]; // @[ToAXI4.scala 243:93]
  wire  d_sel_282 = _d_sel_T_1[282]; // @[ToAXI4.scala 243:93]
  wire  d_sel_283 = _d_sel_T_1[283]; // @[ToAXI4.scala 243:93]
  wire  d_sel_284 = _d_sel_T_1[284]; // @[ToAXI4.scala 243:93]
  wire  d_sel_285 = _d_sel_T_1[285]; // @[ToAXI4.scala 243:93]
  wire  d_sel_286 = _d_sel_T_1[286]; // @[ToAXI4.scala 243:93]
  wire  d_sel_287 = _d_sel_T_1[287]; // @[ToAXI4.scala 243:93]
  wire  d_sel_288 = _d_sel_T_1[288]; // @[ToAXI4.scala 243:93]
  wire  d_sel_289 = _d_sel_T_1[289]; // @[ToAXI4.scala 243:93]
  wire  d_sel_290 = _d_sel_T_1[290]; // @[ToAXI4.scala 243:93]
  wire  d_sel_291 = _d_sel_T_1[291]; // @[ToAXI4.scala 243:93]
  wire  d_sel_292 = _d_sel_T_1[292]; // @[ToAXI4.scala 243:93]
  wire  d_sel_293 = _d_sel_T_1[293]; // @[ToAXI4.scala 243:93]
  wire  d_sel_294 = _d_sel_T_1[294]; // @[ToAXI4.scala 243:93]
  wire  d_sel_295 = _d_sel_T_1[295]; // @[ToAXI4.scala 243:93]
  wire  d_sel_296 = _d_sel_T_1[296]; // @[ToAXI4.scala 243:93]
  wire  d_sel_297 = _d_sel_T_1[297]; // @[ToAXI4.scala 243:93]
  wire  d_sel_298 = _d_sel_T_1[298]; // @[ToAXI4.scala 243:93]
  wire  d_sel_299 = _d_sel_T_1[299]; // @[ToAXI4.scala 243:93]
  wire  d_sel_300 = _d_sel_T_1[300]; // @[ToAXI4.scala 243:93]
  wire  d_sel_301 = _d_sel_T_1[301]; // @[ToAXI4.scala 243:93]
  wire  d_sel_302 = _d_sel_T_1[302]; // @[ToAXI4.scala 243:93]
  wire  d_sel_303 = _d_sel_T_1[303]; // @[ToAXI4.scala 243:93]
  wire  d_sel_304 = _d_sel_T_1[304]; // @[ToAXI4.scala 243:93]
  wire  d_sel_305 = _d_sel_T_1[305]; // @[ToAXI4.scala 243:93]
  wire  d_sel_306 = _d_sel_T_1[306]; // @[ToAXI4.scala 243:93]
  wire  d_sel_307 = _d_sel_T_1[307]; // @[ToAXI4.scala 243:93]
  wire  d_sel_308 = _d_sel_T_1[308]; // @[ToAXI4.scala 243:93]
  wire  d_sel_309 = _d_sel_T_1[309]; // @[ToAXI4.scala 243:93]
  wire  d_sel_310 = _d_sel_T_1[310]; // @[ToAXI4.scala 243:93]
  wire  d_sel_311 = _d_sel_T_1[311]; // @[ToAXI4.scala 243:93]
  wire  d_sel_312 = _d_sel_T_1[312]; // @[ToAXI4.scala 243:93]
  wire  d_sel_313 = _d_sel_T_1[313]; // @[ToAXI4.scala 243:93]
  wire  d_sel_314 = _d_sel_T_1[314]; // @[ToAXI4.scala 243:93]
  wire  d_sel_315 = _d_sel_T_1[315]; // @[ToAXI4.scala 243:93]
  wire  d_sel_316 = _d_sel_T_1[316]; // @[ToAXI4.scala 243:93]
  wire  d_sel_317 = _d_sel_T_1[317]; // @[ToAXI4.scala 243:93]
  wire  d_sel_318 = _d_sel_T_1[318]; // @[ToAXI4.scala 243:93]
  wire  d_sel_319 = _d_sel_T_1[319]; // @[ToAXI4.scala 243:93]
  wire  d_sel_320 = _d_sel_T_1[320]; // @[ToAXI4.scala 243:93]
  wire  d_sel_321 = _d_sel_T_1[321]; // @[ToAXI4.scala 243:93]
  wire  d_sel_322 = _d_sel_T_1[322]; // @[ToAXI4.scala 243:93]
  wire  d_sel_323 = _d_sel_T_1[323]; // @[ToAXI4.scala 243:93]
  wire  d_sel_324 = _d_sel_T_1[324]; // @[ToAXI4.scala 243:93]
  wire  d_sel_325 = _d_sel_T_1[325]; // @[ToAXI4.scala 243:93]
  wire  d_sel_326 = _d_sel_T_1[326]; // @[ToAXI4.scala 243:93]
  wire  d_sel_327 = _d_sel_T_1[327]; // @[ToAXI4.scala 243:93]
  wire  d_sel_328 = _d_sel_T_1[328]; // @[ToAXI4.scala 243:93]
  wire  d_sel_329 = _d_sel_T_1[329]; // @[ToAXI4.scala 243:93]
  wire  d_sel_330 = _d_sel_T_1[330]; // @[ToAXI4.scala 243:93]
  wire  d_sel_331 = _d_sel_T_1[331]; // @[ToAXI4.scala 243:93]
  wire  d_sel_332 = _d_sel_T_1[332]; // @[ToAXI4.scala 243:93]
  wire  d_sel_333 = _d_sel_T_1[333]; // @[ToAXI4.scala 243:93]
  wire  d_sel_334 = _d_sel_T_1[334]; // @[ToAXI4.scala 243:93]
  wire  d_sel_335 = _d_sel_T_1[335]; // @[ToAXI4.scala 243:93]
  wire  d_sel_336 = _d_sel_T_1[336]; // @[ToAXI4.scala 243:93]
  wire  d_sel_337 = _d_sel_T_1[337]; // @[ToAXI4.scala 243:93]
  wire  d_sel_338 = _d_sel_T_1[338]; // @[ToAXI4.scala 243:93]
  wire  d_sel_339 = _d_sel_T_1[339]; // @[ToAXI4.scala 243:93]
  wire  d_sel_340 = _d_sel_T_1[340]; // @[ToAXI4.scala 243:93]
  wire  d_sel_341 = _d_sel_T_1[341]; // @[ToAXI4.scala 243:93]
  wire  d_sel_342 = _d_sel_T_1[342]; // @[ToAXI4.scala 243:93]
  wire  d_sel_343 = _d_sel_T_1[343]; // @[ToAXI4.scala 243:93]
  wire  d_sel_344 = _d_sel_T_1[344]; // @[ToAXI4.scala 243:93]
  wire  d_sel_345 = _d_sel_T_1[345]; // @[ToAXI4.scala 243:93]
  wire  d_sel_346 = _d_sel_T_1[346]; // @[ToAXI4.scala 243:93]
  wire  d_sel_347 = _d_sel_T_1[347]; // @[ToAXI4.scala 243:93]
  wire  d_sel_348 = _d_sel_T_1[348]; // @[ToAXI4.scala 243:93]
  wire  d_sel_349 = _d_sel_T_1[349]; // @[ToAXI4.scala 243:93]
  wire  d_sel_350 = _d_sel_T_1[350]; // @[ToAXI4.scala 243:93]
  wire  d_sel_351 = _d_sel_T_1[351]; // @[ToAXI4.scala 243:93]
  wire  d_sel_352 = _d_sel_T_1[352]; // @[ToAXI4.scala 243:93]
  wire  d_sel_353 = _d_sel_T_1[353]; // @[ToAXI4.scala 243:93]
  wire  d_sel_354 = _d_sel_T_1[354]; // @[ToAXI4.scala 243:93]
  wire  d_sel_355 = _d_sel_T_1[355]; // @[ToAXI4.scala 243:93]
  wire  d_sel_356 = _d_sel_T_1[356]; // @[ToAXI4.scala 243:93]
  wire  d_sel_357 = _d_sel_T_1[357]; // @[ToAXI4.scala 243:93]
  wire  d_sel_358 = _d_sel_T_1[358]; // @[ToAXI4.scala 243:93]
  wire  d_sel_359 = _d_sel_T_1[359]; // @[ToAXI4.scala 243:93]
  wire  d_sel_360 = _d_sel_T_1[360]; // @[ToAXI4.scala 243:93]
  wire  d_sel_361 = _d_sel_T_1[361]; // @[ToAXI4.scala 243:93]
  wire  d_sel_362 = _d_sel_T_1[362]; // @[ToAXI4.scala 243:93]
  wire  d_sel_363 = _d_sel_T_1[363]; // @[ToAXI4.scala 243:93]
  wire  d_sel_364 = _d_sel_T_1[364]; // @[ToAXI4.scala 243:93]
  wire  d_sel_365 = _d_sel_T_1[365]; // @[ToAXI4.scala 243:93]
  wire  d_sel_366 = _d_sel_T_1[366]; // @[ToAXI4.scala 243:93]
  wire  d_sel_367 = _d_sel_T_1[367]; // @[ToAXI4.scala 243:93]
  wire  d_sel_368 = _d_sel_T_1[368]; // @[ToAXI4.scala 243:93]
  wire  d_sel_369 = _d_sel_T_1[369]; // @[ToAXI4.scala 243:93]
  wire  d_sel_370 = _d_sel_T_1[370]; // @[ToAXI4.scala 243:93]
  wire  d_sel_371 = _d_sel_T_1[371]; // @[ToAXI4.scala 243:93]
  wire  d_sel_372 = _d_sel_T_1[372]; // @[ToAXI4.scala 243:93]
  wire  d_sel_373 = _d_sel_T_1[373]; // @[ToAXI4.scala 243:93]
  wire  d_sel_374 = _d_sel_T_1[374]; // @[ToAXI4.scala 243:93]
  wire  d_sel_375 = _d_sel_T_1[375]; // @[ToAXI4.scala 243:93]
  wire  d_sel_376 = _d_sel_T_1[376]; // @[ToAXI4.scala 243:93]
  wire  d_sel_377 = _d_sel_T_1[377]; // @[ToAXI4.scala 243:93]
  wire  d_sel_378 = _d_sel_T_1[378]; // @[ToAXI4.scala 243:93]
  wire  d_sel_379 = _d_sel_T_1[379]; // @[ToAXI4.scala 243:93]
  wire  d_sel_380 = _d_sel_T_1[380]; // @[ToAXI4.scala 243:93]
  wire  d_sel_381 = _d_sel_T_1[381]; // @[ToAXI4.scala 243:93]
  wire  d_sel_382 = _d_sel_T_1[382]; // @[ToAXI4.scala 243:93]
  wire  d_sel_383 = _d_sel_T_1[383]; // @[ToAXI4.scala 243:93]
  wire  d_sel_384 = _d_sel_T_1[384]; // @[ToAXI4.scala 243:93]
  wire  d_sel_385 = _d_sel_T_1[385]; // @[ToAXI4.scala 243:93]
  wire  d_sel_386 = _d_sel_T_1[386]; // @[ToAXI4.scala 243:93]
  wire  d_sel_387 = _d_sel_T_1[387]; // @[ToAXI4.scala 243:93]
  wire  d_sel_388 = _d_sel_T_1[388]; // @[ToAXI4.scala 243:93]
  wire  d_sel_389 = _d_sel_T_1[389]; // @[ToAXI4.scala 243:93]
  wire  d_sel_390 = _d_sel_T_1[390]; // @[ToAXI4.scala 243:93]
  wire  d_sel_391 = _d_sel_T_1[391]; // @[ToAXI4.scala 243:93]
  wire  d_sel_392 = _d_sel_T_1[392]; // @[ToAXI4.scala 243:93]
  wire  d_sel_393 = _d_sel_T_1[393]; // @[ToAXI4.scala 243:93]
  wire  d_sel_394 = _d_sel_T_1[394]; // @[ToAXI4.scala 243:93]
  wire  d_sel_395 = _d_sel_T_1[395]; // @[ToAXI4.scala 243:93]
  wire  d_sel_396 = _d_sel_T_1[396]; // @[ToAXI4.scala 243:93]
  wire  d_sel_397 = _d_sel_T_1[397]; // @[ToAXI4.scala 243:93]
  wire  d_sel_398 = _d_sel_T_1[398]; // @[ToAXI4.scala 243:93]
  wire  d_sel_399 = _d_sel_T_1[399]; // @[ToAXI4.scala 243:93]
  wire  d_sel_400 = _d_sel_T_1[400]; // @[ToAXI4.scala 243:93]
  wire  d_sel_401 = _d_sel_T_1[401]; // @[ToAXI4.scala 243:93]
  wire  d_sel_402 = _d_sel_T_1[402]; // @[ToAXI4.scala 243:93]
  wire  d_sel_403 = _d_sel_T_1[403]; // @[ToAXI4.scala 243:93]
  wire  d_sel_404 = _d_sel_T_1[404]; // @[ToAXI4.scala 243:93]
  wire  d_sel_405 = _d_sel_T_1[405]; // @[ToAXI4.scala 243:93]
  wire  d_sel_406 = _d_sel_T_1[406]; // @[ToAXI4.scala 243:93]
  wire  d_sel_407 = _d_sel_T_1[407]; // @[ToAXI4.scala 243:93]
  wire  d_sel_408 = _d_sel_T_1[408]; // @[ToAXI4.scala 243:93]
  wire  d_sel_409 = _d_sel_T_1[409]; // @[ToAXI4.scala 243:93]
  wire  d_sel_410 = _d_sel_T_1[410]; // @[ToAXI4.scala 243:93]
  wire  d_sel_411 = _d_sel_T_1[411]; // @[ToAXI4.scala 243:93]
  wire  d_sel_412 = _d_sel_T_1[412]; // @[ToAXI4.scala 243:93]
  wire  d_sel_413 = _d_sel_T_1[413]; // @[ToAXI4.scala 243:93]
  wire  d_sel_414 = _d_sel_T_1[414]; // @[ToAXI4.scala 243:93]
  wire  d_sel_415 = _d_sel_T_1[415]; // @[ToAXI4.scala 243:93]
  wire  d_sel_416 = _d_sel_T_1[416]; // @[ToAXI4.scala 243:93]
  wire  d_sel_417 = _d_sel_T_1[417]; // @[ToAXI4.scala 243:93]
  wire  d_sel_418 = _d_sel_T_1[418]; // @[ToAXI4.scala 243:93]
  wire  d_sel_419 = _d_sel_T_1[419]; // @[ToAXI4.scala 243:93]
  wire  d_sel_420 = _d_sel_T_1[420]; // @[ToAXI4.scala 243:93]
  wire  d_sel_421 = _d_sel_T_1[421]; // @[ToAXI4.scala 243:93]
  wire  d_sel_422 = _d_sel_T_1[422]; // @[ToAXI4.scala 243:93]
  wire  d_sel_423 = _d_sel_T_1[423]; // @[ToAXI4.scala 243:93]
  wire  d_sel_424 = _d_sel_T_1[424]; // @[ToAXI4.scala 243:93]
  wire  d_sel_425 = _d_sel_T_1[425]; // @[ToAXI4.scala 243:93]
  wire  d_sel_426 = _d_sel_T_1[426]; // @[ToAXI4.scala 243:93]
  wire  d_sel_427 = _d_sel_T_1[427]; // @[ToAXI4.scala 243:93]
  wire  d_sel_428 = _d_sel_T_1[428]; // @[ToAXI4.scala 243:93]
  wire  d_sel_429 = _d_sel_T_1[429]; // @[ToAXI4.scala 243:93]
  wire  d_sel_430 = _d_sel_T_1[430]; // @[ToAXI4.scala 243:93]
  wire  d_sel_431 = _d_sel_T_1[431]; // @[ToAXI4.scala 243:93]
  wire  d_sel_432 = _d_sel_T_1[432]; // @[ToAXI4.scala 243:93]
  wire  d_sel_433 = _d_sel_T_1[433]; // @[ToAXI4.scala 243:93]
  wire  d_sel_434 = _d_sel_T_1[434]; // @[ToAXI4.scala 243:93]
  wire  d_sel_435 = _d_sel_T_1[435]; // @[ToAXI4.scala 243:93]
  wire  d_sel_436 = _d_sel_T_1[436]; // @[ToAXI4.scala 243:93]
  wire  d_sel_437 = _d_sel_T_1[437]; // @[ToAXI4.scala 243:93]
  wire  d_sel_438 = _d_sel_T_1[438]; // @[ToAXI4.scala 243:93]
  wire  d_sel_439 = _d_sel_T_1[439]; // @[ToAXI4.scala 243:93]
  wire  d_sel_440 = _d_sel_T_1[440]; // @[ToAXI4.scala 243:93]
  wire  d_sel_441 = _d_sel_T_1[441]; // @[ToAXI4.scala 243:93]
  wire  d_sel_442 = _d_sel_T_1[442]; // @[ToAXI4.scala 243:93]
  wire  d_sel_443 = _d_sel_T_1[443]; // @[ToAXI4.scala 243:93]
  wire  d_sel_444 = _d_sel_T_1[444]; // @[ToAXI4.scala 243:93]
  wire  d_sel_445 = _d_sel_T_1[445]; // @[ToAXI4.scala 243:93]
  wire  d_sel_446 = _d_sel_T_1[446]; // @[ToAXI4.scala 243:93]
  wire  d_sel_447 = _d_sel_T_1[447]; // @[ToAXI4.scala 243:93]
  wire  d_sel_448 = _d_sel_T_1[448]; // @[ToAXI4.scala 243:93]
  wire  d_sel_449 = _d_sel_T_1[449]; // @[ToAXI4.scala 243:93]
  wire  d_sel_450 = _d_sel_T_1[450]; // @[ToAXI4.scala 243:93]
  wire  d_sel_451 = _d_sel_T_1[451]; // @[ToAXI4.scala 243:93]
  wire  d_sel_452 = _d_sel_T_1[452]; // @[ToAXI4.scala 243:93]
  wire  d_sel_453 = _d_sel_T_1[453]; // @[ToAXI4.scala 243:93]
  wire  d_sel_454 = _d_sel_T_1[454]; // @[ToAXI4.scala 243:93]
  wire  d_sel_455 = _d_sel_T_1[455]; // @[ToAXI4.scala 243:93]
  wire  d_sel_456 = _d_sel_T_1[456]; // @[ToAXI4.scala 243:93]
  wire  d_sel_457 = _d_sel_T_1[457]; // @[ToAXI4.scala 243:93]
  wire  d_sel_458 = _d_sel_T_1[458]; // @[ToAXI4.scala 243:93]
  wire  d_sel_459 = _d_sel_T_1[459]; // @[ToAXI4.scala 243:93]
  wire  d_sel_460 = _d_sel_T_1[460]; // @[ToAXI4.scala 243:93]
  wire  d_sel_461 = _d_sel_T_1[461]; // @[ToAXI4.scala 243:93]
  wire  d_sel_462 = _d_sel_T_1[462]; // @[ToAXI4.scala 243:93]
  wire  d_sel_463 = _d_sel_T_1[463]; // @[ToAXI4.scala 243:93]
  wire  d_sel_464 = _d_sel_T_1[464]; // @[ToAXI4.scala 243:93]
  wire  d_sel_465 = _d_sel_T_1[465]; // @[ToAXI4.scala 243:93]
  wire  d_sel_466 = _d_sel_T_1[466]; // @[ToAXI4.scala 243:93]
  wire  d_sel_467 = _d_sel_T_1[467]; // @[ToAXI4.scala 243:93]
  wire  d_sel_468 = _d_sel_T_1[468]; // @[ToAXI4.scala 243:93]
  wire  d_sel_469 = _d_sel_T_1[469]; // @[ToAXI4.scala 243:93]
  wire  d_sel_470 = _d_sel_T_1[470]; // @[ToAXI4.scala 243:93]
  wire  d_sel_471 = _d_sel_T_1[471]; // @[ToAXI4.scala 243:93]
  wire  d_sel_472 = _d_sel_T_1[472]; // @[ToAXI4.scala 243:93]
  wire  d_sel_473 = _d_sel_T_1[473]; // @[ToAXI4.scala 243:93]
  wire  d_sel_474 = _d_sel_T_1[474]; // @[ToAXI4.scala 243:93]
  wire  d_sel_475 = _d_sel_T_1[475]; // @[ToAXI4.scala 243:93]
  wire  d_sel_476 = _d_sel_T_1[476]; // @[ToAXI4.scala 243:93]
  wire  d_sel_477 = _d_sel_T_1[477]; // @[ToAXI4.scala 243:93]
  wire  d_sel_478 = _d_sel_T_1[478]; // @[ToAXI4.scala 243:93]
  wire  d_sel_479 = _d_sel_T_1[479]; // @[ToAXI4.scala 243:93]
  wire  d_sel_480 = _d_sel_T_1[480]; // @[ToAXI4.scala 243:93]
  wire  d_sel_481 = _d_sel_T_1[481]; // @[ToAXI4.scala 243:93]
  wire  d_sel_482 = _d_sel_T_1[482]; // @[ToAXI4.scala 243:93]
  wire  d_sel_483 = _d_sel_T_1[483]; // @[ToAXI4.scala 243:93]
  wire  d_sel_484 = _d_sel_T_1[484]; // @[ToAXI4.scala 243:93]
  wire  d_sel_485 = _d_sel_T_1[485]; // @[ToAXI4.scala 243:93]
  wire  d_sel_486 = _d_sel_T_1[486]; // @[ToAXI4.scala 243:93]
  wire  d_sel_487 = _d_sel_T_1[487]; // @[ToAXI4.scala 243:93]
  wire  d_sel_488 = _d_sel_T_1[488]; // @[ToAXI4.scala 243:93]
  wire  d_sel_489 = _d_sel_T_1[489]; // @[ToAXI4.scala 243:93]
  wire  d_sel_490 = _d_sel_T_1[490]; // @[ToAXI4.scala 243:93]
  wire  d_sel_491 = _d_sel_T_1[491]; // @[ToAXI4.scala 243:93]
  wire  d_sel_492 = _d_sel_T_1[492]; // @[ToAXI4.scala 243:93]
  wire  d_sel_493 = _d_sel_T_1[493]; // @[ToAXI4.scala 243:93]
  wire  d_sel_494 = _d_sel_T_1[494]; // @[ToAXI4.scala 243:93]
  wire  d_sel_495 = _d_sel_T_1[495]; // @[ToAXI4.scala 243:93]
  wire  d_sel_496 = _d_sel_T_1[496]; // @[ToAXI4.scala 243:93]
  wire  d_sel_497 = _d_sel_T_1[497]; // @[ToAXI4.scala 243:93]
  wire  d_sel_498 = _d_sel_T_1[498]; // @[ToAXI4.scala 243:93]
  wire  d_sel_499 = _d_sel_T_1[499]; // @[ToAXI4.scala 243:93]
  wire  d_sel_500 = _d_sel_T_1[500]; // @[ToAXI4.scala 243:93]
  wire  d_sel_501 = _d_sel_T_1[501]; // @[ToAXI4.scala 243:93]
  wire  d_sel_502 = _d_sel_T_1[502]; // @[ToAXI4.scala 243:93]
  wire  d_sel_503 = _d_sel_T_1[503]; // @[ToAXI4.scala 243:93]
  wire  d_sel_504 = _d_sel_T_1[504]; // @[ToAXI4.scala 243:93]
  wire  d_sel_505 = _d_sel_T_1[505]; // @[ToAXI4.scala 243:93]
  wire  d_sel_506 = _d_sel_T_1[506]; // @[ToAXI4.scala 243:93]
  wire  d_sel_507 = _d_sel_T_1[507]; // @[ToAXI4.scala 243:93]
  wire  d_sel_508 = _d_sel_T_1[508]; // @[ToAXI4.scala 243:93]
  wire  d_sel_509 = _d_sel_T_1[509]; // @[ToAXI4.scala 243:93]
  wire  d_sel_510 = _d_sel_T_1[510]; // @[ToAXI4.scala 243:93]
  wire  d_sel_511 = _d_sel_T_1[511]; // @[ToAXI4.scala 243:93]
  wire  d_last = r_wins ? auto_out_r_bits_last : 1'h1; // @[ToAXI4.scala 244:23]
  wire  _inc_T = out_arw_ready & out_arw_valid; // @[Decoupled.scala 50:35]
  wire  inc = a_sel_0 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  _dec_T_1 = auto_in_d_ready & bundleIn_0_d_valid; // @[Decoupled.scala 50:35]
  wire  dec = d_sel_0 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  _T_10 = ~reset; // @[ToAXI4.scala 262:16]
  wire  inc_1 = a_sel_1 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_1 = d_sel_1 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_2 = a_sel_2 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_2 = d_sel_2 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_3 = a_sel_3 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_3 = d_sel_3 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_4 = a_sel_4 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_4 = d_sel_4 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_5 = a_sel_5 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_5 = d_sel_5 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_6 = a_sel_6 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_6 = d_sel_6 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_7 = a_sel_7 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_7 = d_sel_7 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_8 = a_sel_8 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_8 = d_sel_8 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_9 = a_sel_9 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_9 = d_sel_9 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_10 = a_sel_10 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_10 = d_sel_10 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_11 = a_sel_11 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_11 = d_sel_11 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_12 = a_sel_12 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_12 = d_sel_12 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_13 = a_sel_13 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_13 = d_sel_13 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_14 = a_sel_14 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_14 = d_sel_14 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_15 = a_sel_15 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_15 = d_sel_15 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_16 = a_sel_16 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_16 = d_sel_16 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_17 = a_sel_17 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_17 = d_sel_17 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_18 = a_sel_18 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_18 = d_sel_18 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_19 = a_sel_19 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_19 = d_sel_19 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_20 = a_sel_20 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_20 = d_sel_20 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_21 = a_sel_21 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_21 = d_sel_21 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_22 = a_sel_22 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_22 = d_sel_22 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_23 = a_sel_23 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_23 = d_sel_23 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_24 = a_sel_24 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_24 = d_sel_24 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_25 = a_sel_25 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_25 = d_sel_25 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_26 = a_sel_26 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_26 = d_sel_26 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_27 = a_sel_27 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_27 = d_sel_27 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_28 = a_sel_28 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_28 = d_sel_28 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_29 = a_sel_29 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_29 = d_sel_29 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_30 = a_sel_30 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_30 = d_sel_30 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_31 = a_sel_31 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_31 = d_sel_31 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_32 = a_sel_32 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_32 = d_sel_32 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_33 = a_sel_33 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_33 = d_sel_33 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_34 = a_sel_34 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_34 = d_sel_34 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_35 = a_sel_35 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_35 = d_sel_35 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_36 = a_sel_36 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_36 = d_sel_36 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_37 = a_sel_37 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_37 = d_sel_37 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_38 = a_sel_38 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_38 = d_sel_38 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_39 = a_sel_39 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_39 = d_sel_39 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_40 = a_sel_40 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_40 = d_sel_40 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_41 = a_sel_41 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_41 = d_sel_41 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_42 = a_sel_42 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_42 = d_sel_42 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_43 = a_sel_43 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_43 = d_sel_43 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_44 = a_sel_44 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_44 = d_sel_44 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_45 = a_sel_45 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_45 = d_sel_45 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_46 = a_sel_46 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_46 = d_sel_46 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_47 = a_sel_47 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_47 = d_sel_47 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_48 = a_sel_48 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_48 = d_sel_48 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_49 = a_sel_49 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_49 = d_sel_49 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_50 = a_sel_50 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_50 = d_sel_50 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_51 = a_sel_51 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_51 = d_sel_51 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_52 = a_sel_52 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_52 = d_sel_52 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_53 = a_sel_53 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_53 = d_sel_53 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_54 = a_sel_54 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_54 = d_sel_54 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_55 = a_sel_55 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_55 = d_sel_55 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_56 = a_sel_56 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_56 = d_sel_56 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_57 = a_sel_57 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_57 = d_sel_57 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_58 = a_sel_58 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_58 = d_sel_58 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_59 = a_sel_59 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_59 = d_sel_59 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_60 = a_sel_60 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_60 = d_sel_60 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_61 = a_sel_61 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_61 = d_sel_61 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_62 = a_sel_62 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_62 = d_sel_62 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_63 = a_sel_63 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_63 = d_sel_63 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_64 = a_sel_64 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_64 = d_sel_64 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_65 = a_sel_65 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_65 = d_sel_65 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_66 = a_sel_66 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_66 = d_sel_66 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_67 = a_sel_67 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_67 = d_sel_67 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_68 = a_sel_68 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_68 = d_sel_68 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_69 = a_sel_69 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_69 = d_sel_69 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_70 = a_sel_70 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_70 = d_sel_70 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_71 = a_sel_71 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_71 = d_sel_71 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_72 = a_sel_72 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_72 = d_sel_72 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_73 = a_sel_73 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_73 = d_sel_73 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_74 = a_sel_74 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_74 = d_sel_74 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_75 = a_sel_75 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_75 = d_sel_75 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_76 = a_sel_76 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_76 = d_sel_76 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_77 = a_sel_77 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_77 = d_sel_77 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_78 = a_sel_78 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_78 = d_sel_78 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_79 = a_sel_79 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_79 = d_sel_79 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_80 = a_sel_80 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_80 = d_sel_80 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_81 = a_sel_81 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_81 = d_sel_81 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_82 = a_sel_82 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_82 = d_sel_82 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_83 = a_sel_83 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_83 = d_sel_83 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_84 = a_sel_84 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_84 = d_sel_84 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_85 = a_sel_85 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_85 = d_sel_85 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_86 = a_sel_86 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_86 = d_sel_86 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_87 = a_sel_87 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_87 = d_sel_87 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_88 = a_sel_88 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_88 = d_sel_88 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_89 = a_sel_89 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_89 = d_sel_89 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_90 = a_sel_90 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_90 = d_sel_90 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_91 = a_sel_91 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_91 = d_sel_91 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_92 = a_sel_92 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_92 = d_sel_92 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_93 = a_sel_93 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_93 = d_sel_93 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_94 = a_sel_94 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_94 = d_sel_94 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_95 = a_sel_95 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_95 = d_sel_95 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_96 = a_sel_96 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_96 = d_sel_96 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_97 = a_sel_97 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_97 = d_sel_97 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_98 = a_sel_98 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_98 = d_sel_98 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_99 = a_sel_99 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_99 = d_sel_99 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_100 = a_sel_100 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_100 = d_sel_100 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_101 = a_sel_101 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_101 = d_sel_101 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_102 = a_sel_102 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_102 = d_sel_102 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_103 = a_sel_103 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_103 = d_sel_103 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_104 = a_sel_104 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_104 = d_sel_104 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_105 = a_sel_105 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_105 = d_sel_105 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_106 = a_sel_106 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_106 = d_sel_106 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_107 = a_sel_107 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_107 = d_sel_107 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_108 = a_sel_108 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_108 = d_sel_108 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_109 = a_sel_109 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_109 = d_sel_109 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_110 = a_sel_110 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_110 = d_sel_110 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_111 = a_sel_111 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_111 = d_sel_111 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_112 = a_sel_112 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_112 = d_sel_112 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_113 = a_sel_113 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_113 = d_sel_113 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_114 = a_sel_114 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_114 = d_sel_114 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_115 = a_sel_115 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_115 = d_sel_115 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_116 = a_sel_116 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_116 = d_sel_116 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_117 = a_sel_117 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_117 = d_sel_117 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_118 = a_sel_118 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_118 = d_sel_118 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_119 = a_sel_119 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_119 = d_sel_119 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_120 = a_sel_120 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_120 = d_sel_120 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_121 = a_sel_121 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_121 = d_sel_121 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_122 = a_sel_122 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_122 = d_sel_122 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_123 = a_sel_123 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_123 = d_sel_123 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_124 = a_sel_124 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_124 = d_sel_124 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_125 = a_sel_125 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_125 = d_sel_125 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_126 = a_sel_126 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_126 = d_sel_126 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_127 = a_sel_127 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_127 = d_sel_127 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_128 = a_sel_128 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_128 = d_sel_128 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_129 = a_sel_129 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_129 = d_sel_129 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_130 = a_sel_130 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_130 = d_sel_130 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_131 = a_sel_131 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_131 = d_sel_131 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_132 = a_sel_132 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_132 = d_sel_132 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_133 = a_sel_133 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_133 = d_sel_133 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_134 = a_sel_134 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_134 = d_sel_134 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_135 = a_sel_135 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_135 = d_sel_135 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_136 = a_sel_136 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_136 = d_sel_136 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_137 = a_sel_137 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_137 = d_sel_137 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_138 = a_sel_138 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_138 = d_sel_138 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_139 = a_sel_139 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_139 = d_sel_139 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_140 = a_sel_140 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_140 = d_sel_140 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_141 = a_sel_141 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_141 = d_sel_141 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_142 = a_sel_142 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_142 = d_sel_142 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_143 = a_sel_143 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_143 = d_sel_143 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_144 = a_sel_144 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_144 = d_sel_144 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_145 = a_sel_145 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_145 = d_sel_145 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_146 = a_sel_146 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_146 = d_sel_146 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_147 = a_sel_147 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_147 = d_sel_147 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_148 = a_sel_148 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_148 = d_sel_148 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_149 = a_sel_149 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_149 = d_sel_149 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_150 = a_sel_150 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_150 = d_sel_150 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_151 = a_sel_151 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_151 = d_sel_151 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_152 = a_sel_152 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_152 = d_sel_152 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_153 = a_sel_153 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_153 = d_sel_153 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_154 = a_sel_154 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_154 = d_sel_154 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_155 = a_sel_155 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_155 = d_sel_155 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_156 = a_sel_156 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_156 = d_sel_156 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_157 = a_sel_157 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_157 = d_sel_157 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_158 = a_sel_158 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_158 = d_sel_158 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_159 = a_sel_159 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_159 = d_sel_159 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_160 = a_sel_160 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_160 = d_sel_160 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_161 = a_sel_161 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_161 = d_sel_161 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_162 = a_sel_162 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_162 = d_sel_162 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_163 = a_sel_163 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_163 = d_sel_163 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_164 = a_sel_164 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_164 = d_sel_164 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_165 = a_sel_165 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_165 = d_sel_165 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_166 = a_sel_166 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_166 = d_sel_166 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_167 = a_sel_167 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_167 = d_sel_167 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_168 = a_sel_168 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_168 = d_sel_168 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_169 = a_sel_169 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_169 = d_sel_169 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_170 = a_sel_170 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_170 = d_sel_170 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_171 = a_sel_171 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_171 = d_sel_171 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_172 = a_sel_172 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_172 = d_sel_172 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_173 = a_sel_173 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_173 = d_sel_173 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_174 = a_sel_174 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_174 = d_sel_174 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_175 = a_sel_175 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_175 = d_sel_175 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_176 = a_sel_176 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_176 = d_sel_176 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_177 = a_sel_177 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_177 = d_sel_177 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_178 = a_sel_178 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_178 = d_sel_178 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_179 = a_sel_179 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_179 = d_sel_179 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_180 = a_sel_180 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_180 = d_sel_180 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_181 = a_sel_181 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_181 = d_sel_181 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_182 = a_sel_182 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_182 = d_sel_182 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_183 = a_sel_183 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_183 = d_sel_183 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_184 = a_sel_184 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_184 = d_sel_184 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_185 = a_sel_185 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_185 = d_sel_185 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_186 = a_sel_186 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_186 = d_sel_186 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_187 = a_sel_187 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_187 = d_sel_187 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_188 = a_sel_188 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_188 = d_sel_188 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_189 = a_sel_189 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_189 = d_sel_189 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_190 = a_sel_190 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_190 = d_sel_190 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_191 = a_sel_191 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_191 = d_sel_191 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_192 = a_sel_192 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_192 = d_sel_192 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_193 = a_sel_193 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_193 = d_sel_193 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_194 = a_sel_194 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_194 = d_sel_194 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_195 = a_sel_195 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_195 = d_sel_195 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_196 = a_sel_196 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_196 = d_sel_196 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_197 = a_sel_197 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_197 = d_sel_197 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_198 = a_sel_198 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_198 = d_sel_198 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_199 = a_sel_199 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_199 = d_sel_199 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_200 = a_sel_200 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_200 = d_sel_200 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_201 = a_sel_201 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_201 = d_sel_201 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_202 = a_sel_202 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_202 = d_sel_202 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_203 = a_sel_203 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_203 = d_sel_203 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_204 = a_sel_204 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_204 = d_sel_204 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_205 = a_sel_205 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_205 = d_sel_205 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_206 = a_sel_206 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_206 = d_sel_206 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_207 = a_sel_207 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_207 = d_sel_207 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_208 = a_sel_208 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_208 = d_sel_208 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_209 = a_sel_209 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_209 = d_sel_209 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_210 = a_sel_210 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_210 = d_sel_210 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_211 = a_sel_211 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_211 = d_sel_211 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_212 = a_sel_212 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_212 = d_sel_212 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_213 = a_sel_213 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_213 = d_sel_213 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_214 = a_sel_214 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_214 = d_sel_214 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_215 = a_sel_215 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_215 = d_sel_215 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_216 = a_sel_216 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_216 = d_sel_216 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_217 = a_sel_217 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_217 = d_sel_217 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_218 = a_sel_218 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_218 = d_sel_218 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_219 = a_sel_219 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_219 = d_sel_219 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_220 = a_sel_220 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_220 = d_sel_220 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_221 = a_sel_221 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_221 = d_sel_221 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_222 = a_sel_222 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_222 = d_sel_222 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_223 = a_sel_223 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_223 = d_sel_223 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_224 = a_sel_224 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_224 = d_sel_224 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_225 = a_sel_225 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_225 = d_sel_225 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_226 = a_sel_226 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_226 = d_sel_226 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_227 = a_sel_227 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_227 = d_sel_227 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_228 = a_sel_228 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_228 = d_sel_228 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_229 = a_sel_229 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_229 = d_sel_229 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_230 = a_sel_230 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_230 = d_sel_230 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_231 = a_sel_231 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_231 = d_sel_231 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_232 = a_sel_232 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_232 = d_sel_232 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_233 = a_sel_233 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_233 = d_sel_233 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_234 = a_sel_234 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_234 = d_sel_234 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_235 = a_sel_235 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_235 = d_sel_235 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_236 = a_sel_236 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_236 = d_sel_236 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_237 = a_sel_237 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_237 = d_sel_237 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_238 = a_sel_238 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_238 = d_sel_238 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_239 = a_sel_239 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_239 = d_sel_239 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_240 = a_sel_240 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_240 = d_sel_240 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_241 = a_sel_241 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_241 = d_sel_241 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_242 = a_sel_242 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_242 = d_sel_242 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_243 = a_sel_243 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_243 = d_sel_243 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_244 = a_sel_244 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_244 = d_sel_244 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_245 = a_sel_245 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_245 = d_sel_245 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_246 = a_sel_246 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_246 = d_sel_246 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_247 = a_sel_247 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_247 = d_sel_247 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_248 = a_sel_248 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_248 = d_sel_248 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_249 = a_sel_249 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_249 = d_sel_249 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_250 = a_sel_250 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_250 = d_sel_250 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_251 = a_sel_251 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_251 = d_sel_251 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_252 = a_sel_252 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_252 = d_sel_252 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_253 = a_sel_253 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_253 = d_sel_253 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_254 = a_sel_254 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_254 = d_sel_254 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_255 = a_sel_255 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_255 = d_sel_255 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_256 = a_sel_256 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_256 = d_sel_256 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_257 = a_sel_257 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_257 = d_sel_257 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_258 = a_sel_258 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_258 = d_sel_258 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_259 = a_sel_259 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_259 = d_sel_259 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_260 = a_sel_260 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_260 = d_sel_260 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_261 = a_sel_261 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_261 = d_sel_261 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_262 = a_sel_262 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_262 = d_sel_262 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_263 = a_sel_263 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_263 = d_sel_263 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_264 = a_sel_264 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_264 = d_sel_264 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_265 = a_sel_265 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_265 = d_sel_265 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_266 = a_sel_266 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_266 = d_sel_266 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_267 = a_sel_267 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_267 = d_sel_267 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_268 = a_sel_268 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_268 = d_sel_268 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_269 = a_sel_269 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_269 = d_sel_269 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_270 = a_sel_270 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_270 = d_sel_270 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_271 = a_sel_271 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_271 = d_sel_271 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_272 = a_sel_272 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_272 = d_sel_272 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_273 = a_sel_273 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_273 = d_sel_273 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_274 = a_sel_274 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_274 = d_sel_274 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_275 = a_sel_275 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_275 = d_sel_275 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_276 = a_sel_276 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_276 = d_sel_276 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_277 = a_sel_277 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_277 = d_sel_277 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_278 = a_sel_278 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_278 = d_sel_278 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_279 = a_sel_279 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_279 = d_sel_279 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_280 = a_sel_280 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_280 = d_sel_280 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_281 = a_sel_281 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_281 = d_sel_281 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_282 = a_sel_282 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_282 = d_sel_282 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_283 = a_sel_283 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_283 = d_sel_283 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_284 = a_sel_284 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_284 = d_sel_284 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_285 = a_sel_285 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_285 = d_sel_285 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_286 = a_sel_286 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_286 = d_sel_286 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_287 = a_sel_287 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_287 = d_sel_287 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_288 = a_sel_288 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_288 = d_sel_288 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_289 = a_sel_289 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_289 = d_sel_289 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_290 = a_sel_290 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_290 = d_sel_290 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_291 = a_sel_291 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_291 = d_sel_291 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_292 = a_sel_292 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_292 = d_sel_292 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_293 = a_sel_293 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_293 = d_sel_293 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_294 = a_sel_294 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_294 = d_sel_294 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_295 = a_sel_295 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_295 = d_sel_295 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_296 = a_sel_296 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_296 = d_sel_296 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_297 = a_sel_297 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_297 = d_sel_297 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_298 = a_sel_298 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_298 = d_sel_298 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_299 = a_sel_299 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_299 = d_sel_299 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_300 = a_sel_300 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_300 = d_sel_300 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_301 = a_sel_301 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_301 = d_sel_301 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_302 = a_sel_302 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_302 = d_sel_302 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_303 = a_sel_303 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_303 = d_sel_303 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_304 = a_sel_304 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_304 = d_sel_304 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_305 = a_sel_305 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_305 = d_sel_305 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_306 = a_sel_306 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_306 = d_sel_306 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_307 = a_sel_307 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_307 = d_sel_307 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_308 = a_sel_308 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_308 = d_sel_308 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_309 = a_sel_309 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_309 = d_sel_309 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_310 = a_sel_310 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_310 = d_sel_310 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_311 = a_sel_311 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_311 = d_sel_311 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_312 = a_sel_312 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_312 = d_sel_312 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_313 = a_sel_313 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_313 = d_sel_313 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_314 = a_sel_314 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_314 = d_sel_314 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_315 = a_sel_315 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_315 = d_sel_315 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_316 = a_sel_316 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_316 = d_sel_316 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_317 = a_sel_317 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_317 = d_sel_317 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_318 = a_sel_318 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_318 = d_sel_318 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_319 = a_sel_319 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_319 = d_sel_319 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_320 = a_sel_320 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_320 = d_sel_320 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_321 = a_sel_321 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_321 = d_sel_321 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_322 = a_sel_322 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_322 = d_sel_322 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_323 = a_sel_323 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_323 = d_sel_323 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_324 = a_sel_324 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_324 = d_sel_324 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_325 = a_sel_325 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_325 = d_sel_325 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_326 = a_sel_326 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_326 = d_sel_326 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_327 = a_sel_327 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_327 = d_sel_327 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_328 = a_sel_328 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_328 = d_sel_328 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_329 = a_sel_329 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_329 = d_sel_329 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_330 = a_sel_330 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_330 = d_sel_330 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_331 = a_sel_331 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_331 = d_sel_331 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_332 = a_sel_332 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_332 = d_sel_332 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_333 = a_sel_333 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_333 = d_sel_333 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_334 = a_sel_334 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_334 = d_sel_334 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_335 = a_sel_335 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_335 = d_sel_335 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_336 = a_sel_336 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_336 = d_sel_336 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_337 = a_sel_337 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_337 = d_sel_337 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_338 = a_sel_338 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_338 = d_sel_338 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_339 = a_sel_339 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_339 = d_sel_339 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_340 = a_sel_340 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_340 = d_sel_340 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_341 = a_sel_341 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_341 = d_sel_341 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_342 = a_sel_342 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_342 = d_sel_342 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_343 = a_sel_343 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_343 = d_sel_343 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_344 = a_sel_344 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_344 = d_sel_344 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_345 = a_sel_345 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_345 = d_sel_345 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_346 = a_sel_346 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_346 = d_sel_346 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_347 = a_sel_347 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_347 = d_sel_347 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_348 = a_sel_348 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_348 = d_sel_348 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_349 = a_sel_349 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_349 = d_sel_349 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_350 = a_sel_350 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_350 = d_sel_350 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_351 = a_sel_351 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_351 = d_sel_351 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_352 = a_sel_352 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_352 = d_sel_352 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_353 = a_sel_353 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_353 = d_sel_353 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_354 = a_sel_354 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_354 = d_sel_354 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_355 = a_sel_355 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_355 = d_sel_355 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_356 = a_sel_356 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_356 = d_sel_356 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_357 = a_sel_357 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_357 = d_sel_357 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_358 = a_sel_358 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_358 = d_sel_358 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_359 = a_sel_359 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_359 = d_sel_359 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_360 = a_sel_360 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_360 = d_sel_360 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_361 = a_sel_361 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_361 = d_sel_361 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_362 = a_sel_362 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_362 = d_sel_362 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_363 = a_sel_363 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_363 = d_sel_363 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_364 = a_sel_364 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_364 = d_sel_364 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_365 = a_sel_365 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_365 = d_sel_365 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_366 = a_sel_366 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_366 = d_sel_366 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_367 = a_sel_367 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_367 = d_sel_367 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_368 = a_sel_368 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_368 = d_sel_368 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_369 = a_sel_369 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_369 = d_sel_369 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_370 = a_sel_370 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_370 = d_sel_370 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_371 = a_sel_371 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_371 = d_sel_371 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_372 = a_sel_372 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_372 = d_sel_372 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_373 = a_sel_373 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_373 = d_sel_373 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_374 = a_sel_374 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_374 = d_sel_374 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_375 = a_sel_375 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_375 = d_sel_375 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_376 = a_sel_376 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_376 = d_sel_376 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_377 = a_sel_377 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_377 = d_sel_377 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_378 = a_sel_378 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_378 = d_sel_378 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_379 = a_sel_379 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_379 = d_sel_379 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_380 = a_sel_380 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_380 = d_sel_380 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_381 = a_sel_381 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_381 = d_sel_381 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_382 = a_sel_382 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_382 = d_sel_382 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_383 = a_sel_383 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_383 = d_sel_383 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_384 = a_sel_384 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_384 = d_sel_384 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_385 = a_sel_385 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_385 = d_sel_385 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_386 = a_sel_386 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_386 = d_sel_386 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_387 = a_sel_387 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_387 = d_sel_387 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_388 = a_sel_388 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_388 = d_sel_388 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_389 = a_sel_389 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_389 = d_sel_389 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_390 = a_sel_390 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_390 = d_sel_390 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_391 = a_sel_391 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_391 = d_sel_391 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_392 = a_sel_392 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_392 = d_sel_392 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_393 = a_sel_393 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_393 = d_sel_393 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_394 = a_sel_394 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_394 = d_sel_394 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_395 = a_sel_395 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_395 = d_sel_395 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_396 = a_sel_396 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_396 = d_sel_396 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_397 = a_sel_397 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_397 = d_sel_397 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_398 = a_sel_398 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_398 = d_sel_398 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_399 = a_sel_399 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_399 = d_sel_399 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_400 = a_sel_400 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_400 = d_sel_400 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_401 = a_sel_401 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_401 = d_sel_401 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_402 = a_sel_402 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_402 = d_sel_402 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_403 = a_sel_403 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_403 = d_sel_403 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_404 = a_sel_404 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_404 = d_sel_404 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_405 = a_sel_405 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_405 = d_sel_405 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_406 = a_sel_406 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_406 = d_sel_406 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_407 = a_sel_407 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_407 = d_sel_407 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_408 = a_sel_408 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_408 = d_sel_408 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_409 = a_sel_409 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_409 = d_sel_409 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_410 = a_sel_410 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_410 = d_sel_410 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_411 = a_sel_411 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_411 = d_sel_411 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_412 = a_sel_412 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_412 = d_sel_412 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_413 = a_sel_413 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_413 = d_sel_413 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_414 = a_sel_414 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_414 = d_sel_414 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_415 = a_sel_415 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_415 = d_sel_415 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_416 = a_sel_416 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_416 = d_sel_416 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_417 = a_sel_417 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_417 = d_sel_417 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_418 = a_sel_418 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_418 = d_sel_418 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_419 = a_sel_419 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_419 = d_sel_419 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_420 = a_sel_420 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_420 = d_sel_420 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_421 = a_sel_421 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_421 = d_sel_421 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_422 = a_sel_422 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_422 = d_sel_422 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_423 = a_sel_423 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_423 = d_sel_423 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_424 = a_sel_424 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_424 = d_sel_424 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_425 = a_sel_425 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_425 = d_sel_425 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_426 = a_sel_426 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_426 = d_sel_426 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_427 = a_sel_427 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_427 = d_sel_427 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_428 = a_sel_428 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_428 = d_sel_428 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_429 = a_sel_429 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_429 = d_sel_429 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_430 = a_sel_430 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_430 = d_sel_430 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_431 = a_sel_431 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_431 = d_sel_431 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_432 = a_sel_432 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_432 = d_sel_432 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_433 = a_sel_433 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_433 = d_sel_433 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_434 = a_sel_434 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_434 = d_sel_434 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_435 = a_sel_435 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_435 = d_sel_435 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_436 = a_sel_436 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_436 = d_sel_436 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_437 = a_sel_437 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_437 = d_sel_437 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_438 = a_sel_438 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_438 = d_sel_438 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_439 = a_sel_439 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_439 = d_sel_439 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_440 = a_sel_440 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_440 = d_sel_440 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_441 = a_sel_441 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_441 = d_sel_441 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_442 = a_sel_442 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_442 = d_sel_442 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_443 = a_sel_443 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_443 = d_sel_443 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_444 = a_sel_444 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_444 = d_sel_444 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_445 = a_sel_445 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_445 = d_sel_445 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_446 = a_sel_446 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_446 = d_sel_446 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_447 = a_sel_447 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_447 = d_sel_447 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_448 = a_sel_448 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_448 = d_sel_448 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_449 = a_sel_449 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_449 = d_sel_449 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_450 = a_sel_450 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_450 = d_sel_450 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_451 = a_sel_451 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_451 = d_sel_451 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_452 = a_sel_452 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_452 = d_sel_452 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_453 = a_sel_453 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_453 = d_sel_453 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_454 = a_sel_454 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_454 = d_sel_454 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_455 = a_sel_455 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_455 = d_sel_455 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_456 = a_sel_456 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_456 = d_sel_456 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_457 = a_sel_457 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_457 = d_sel_457 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_458 = a_sel_458 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_458 = d_sel_458 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_459 = a_sel_459 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_459 = d_sel_459 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_460 = a_sel_460 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_460 = d_sel_460 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_461 = a_sel_461 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_461 = d_sel_461 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_462 = a_sel_462 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_462 = d_sel_462 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_463 = a_sel_463 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_463 = d_sel_463 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_464 = a_sel_464 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_464 = d_sel_464 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_465 = a_sel_465 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_465 = d_sel_465 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_466 = a_sel_466 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_466 = d_sel_466 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_467 = a_sel_467 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_467 = d_sel_467 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_468 = a_sel_468 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_468 = d_sel_468 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_469 = a_sel_469 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_469 = d_sel_469 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_470 = a_sel_470 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_470 = d_sel_470 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_471 = a_sel_471 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_471 = d_sel_471 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_472 = a_sel_472 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_472 = d_sel_472 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_473 = a_sel_473 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_473 = d_sel_473 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_474 = a_sel_474 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_474 = d_sel_474 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_475 = a_sel_475 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_475 = d_sel_475 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_476 = a_sel_476 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_476 = d_sel_476 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_477 = a_sel_477 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_477 = d_sel_477 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_478 = a_sel_478 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_478 = d_sel_478 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_479 = a_sel_479 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_479 = d_sel_479 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_480 = a_sel_480 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_480 = d_sel_480 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_481 = a_sel_481 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_481 = d_sel_481 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_482 = a_sel_482 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_482 = d_sel_482 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_483 = a_sel_483 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_483 = d_sel_483 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_484 = a_sel_484 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_484 = d_sel_484 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_485 = a_sel_485 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_485 = d_sel_485 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_486 = a_sel_486 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_486 = d_sel_486 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_487 = a_sel_487 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_487 = d_sel_487 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_488 = a_sel_488 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_488 = d_sel_488 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_489 = a_sel_489 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_489 = d_sel_489 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_490 = a_sel_490 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_490 = d_sel_490 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_491 = a_sel_491 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_491 = d_sel_491 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_492 = a_sel_492 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_492 = d_sel_492 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_493 = a_sel_493 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_493 = d_sel_493 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_494 = a_sel_494 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_494 = d_sel_494 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_495 = a_sel_495 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_495 = d_sel_495 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_496 = a_sel_496 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_496 = d_sel_496 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_497 = a_sel_497 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_497 = d_sel_497 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_498 = a_sel_498 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_498 = d_sel_498 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_499 = a_sel_499 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_499 = d_sel_499 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_500 = a_sel_500 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_500 = d_sel_500 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_501 = a_sel_501 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_501 = d_sel_501 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_502 = a_sel_502 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_502 = d_sel_502 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_503 = a_sel_503 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_503 = d_sel_503 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_504 = a_sel_504 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_504 = d_sel_504 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_505 = a_sel_505 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_505 = d_sel_505 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_506 = a_sel_506 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_506 = d_sel_506 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_507 = a_sel_507 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_507 = d_sel_507 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_508 = a_sel_508 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_508 = d_sel_508 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_509 = a_sel_509 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_509 = d_sel_509 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_510 = a_sel_510 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_510 = d_sel_510 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  wire  inc_511 = a_sel_511 & _inc_T; // @[ToAXI4.scala 258:22]
  wire  dec_511 = d_sel_511 & d_last & _dec_T_1; // @[ToAXI4.scala 259:32]
  reg [19:0] TLToAXI4_covState; // @[Register tracking TLToAXI4 state]
  reg  TLToAXI4_covMap [0:1048575]; // @[Coverage map for TLToAXI4]
  wire  TLToAXI4_covMap_read_en; // @[Coverage map for TLToAXI4]
  wire [19:0] TLToAXI4_covMap_read_addr; // @[Coverage map for TLToAXI4]
  wire  TLToAXI4_covMap_read_data; // @[Coverage map for TLToAXI4]
  wire  TLToAXI4_covMap_write_data; // @[Coverage map for TLToAXI4]
  wire [19:0] TLToAXI4_covMap_write_addr; // @[Coverage map for TLToAXI4]
  wire  TLToAXI4_covMap_write_mask; // @[Coverage map for TLToAXI4]
  wire  TLToAXI4_covMap_write_en; // @[Coverage map for TLToAXI4]
  reg [29:0] TLToAXI4_covSum; // @[Sum of coverage map]
  wire [10:0] count_331_shl;
  wire [19:0] count_331_pad;
  wire [17:0] count_401_shl;
  wire [19:0] count_401_pad;
  wire [18:0] count_227_shl;
  wire [19:0] count_227_pad;
  wire [2:0] count_383_shl;
  wire [19:0] count_383_pad;
  wire [7:0] count_195_shl;
  wire [19:0] count_195_pad;
  wire [18:0] count_417_shl;
  wire [19:0] count_417_pad;
  wire [10:0] count_121_shl;
  wire [19:0] count_121_pad;
  wire [12:0] count_447_shl;
  wire [19:0] count_447_pad;
  wire [12:0] count_482_shl;
  wire [19:0] count_482_pad;
  wire  count_26_shl;
  wire [19:0] count_26_pad;
  wire [17:0] count_391_shl;
  wire [19:0] count_391_pad;
  wire [18:0] count_284_shl;
  wire [19:0] count_284_pad;
  wire [4:0] count_204_shl;
  wire [19:0] count_204_pad;
  wire [13:0] count_199_shl;
  wire [19:0] count_199_pad;
  wire [4:0] count_373_shl;
  wire [19:0] count_373_pad;
  wire [9:0] count_394_shl;
  wire [19:0] count_394_pad;
  wire [13:0] count_411_shl;
  wire [19:0] count_411_pad;
  wire [16:0] count_120_shl;
  wire [19:0] count_120_pad;
  wire [17:0] count_503_shl;
  wire [19:0] count_503_pad;
  wire [3:0] count_70_shl;
  wire [19:0] count_70_pad;
  wire [8:0] count_270_shl;
  wire [19:0] count_270_pad;
  wire [14:0] count_372_shl;
  wire [19:0] count_372_pad;
  wire [12:0] count_474_shl;
  wire [19:0] count_474_pad;
  wire [17:0] count_421_shl;
  wire [19:0] count_421_pad;
  wire [6:0] count_501_shl;
  wire [19:0] count_501_pad;
  wire [2:0] count_154_shl;
  wire [19:0] count_154_pad;
  wire [9:0] count_329_shl;
  wire [19:0] count_329_pad;
  wire [3:0] count_117_shl;
  wire [19:0] count_117_pad;
  wire [12:0] count_297_shl;
  wire [19:0] count_297_pad;
  wire [4:0] count_202_shl;
  wire [19:0] count_202_pad;
  wire [5:0] count_50_shl;
  wire [19:0] count_50_pad;
  wire [11:0] count_184_shl;
  wire [19:0] count_184_pad;
  wire [7:0] count_263_shl;
  wire [19:0] count_263_pad;
  wire [19:0] count_313_shl;
  wire [19:0] count_313_pad;
  wire [12:0] count_168_shl;
  wire [19:0] count_168_pad;
  wire [2:0] count_305_shl;
  wire [19:0] count_305_pad;
  wire [1:0] count_38_shl;
  wire [19:0] count_38_pad;
  wire [1:0] count_310_shl;
  wire [19:0] count_310_pad;
  wire [16:0] count_317_shl;
  wire [19:0] count_317_pad;
  wire  count_393_shl;
  wire [19:0] count_393_pad;
  wire [8:0] count_182_shl;
  wire [19:0] count_182_pad;
  wire [12:0] count_357_shl;
  wire [19:0] count_357_pad;
  wire [15:0] count_423_shl;
  wire [19:0] count_423_pad;
  wire [19:0] count_37_shl;
  wire [19:0] count_37_pad;
  wire [4:0] count_31_shl;
  wire [19:0] count_31_pad;
  wire [6:0] count_61_shl;
  wire [19:0] count_61_pad;
  wire [15:0] count_333_shl;
  wire [19:0] count_333_pad;
  wire  count_296_shl;
  wire [19:0] count_296_pad;
  wire [13:0] count_222_shl;
  wire [19:0] count_222_pad;
  wire [17:0] count_477_shl;
  wire [19:0] count_477_pad;
  wire [14:0] count_498_shl;
  wire [19:0] count_498_pad;
  wire [10:0] count_422_shl;
  wire [19:0] count_422_pad;
  wire [3:0] count_67_shl;
  wire [19:0] count_67_pad;
  wire [1:0] count_420_shl;
  wire [19:0] count_420_pad;
  wire [2:0] count_293_shl;
  wire [19:0] count_293_pad;
  wire [15:0] count_242_shl;
  wire [19:0] count_242_pad;
  wire [1:0] count_64_shl;
  wire [19:0] count_64_pad;
  wire [7:0] count_223_shl;
  wire [19:0] count_223_pad;
  wire [19:0] count_352_shl;
  wire [19:0] count_352_pad;
  wire [9:0] count_153_shl;
  wire [19:0] count_153_pad;
  wire [14:0] count_118_shl;
  wire [19:0] count_118_pad;
  wire [1:0] count_139_shl;
  wire [19:0] count_139_pad;
  wire [8:0] count_467_shl;
  wire [19:0] count_467_pad;
  wire [2:0] count_386_shl;
  wire [19:0] count_386_pad;
  wire [6:0] count_434_shl;
  wire [19:0] count_434_pad;
  wire [16:0] count_51_shl;
  wire [19:0] count_51_pad;
  wire [13:0] count_129_shl;
  wire [19:0] count_129_pad;
  wire [5:0] count_378_shl;
  wire [19:0] count_378_pad;
  wire [10:0] count_186_shl;
  wire [19:0] count_186_pad;
  wire [9:0] count_101_shl;
  wire [19:0] count_101_pad;
  wire [19:0] count_229_shl;
  wire [19:0] count_229_pad;
  wire [10:0] count_280_shl;
  wire [19:0] count_280_pad;
  wire [11:0] count_403_shl;
  wire [19:0] count_403_pad;
  wire [8:0] count_330_shl;
  wire [19:0] count_330_pad;
  wire [10:0] count_398_shl;
  wire [19:0] count_398_pad;
  wire [4:0] count_307_shl;
  wire [19:0] count_307_pad;
  wire [1:0] count_216_shl;
  wire [19:0] count_216_pad;
  wire [6:0] count_400_shl;
  wire [19:0] count_400_pad;
  wire [3:0] count_304_shl;
  wire [19:0] count_304_pad;
  wire [13:0] count_131_shl;
  wire [19:0] count_131_pad;
  wire [9:0] count_282_shl;
  wire [19:0] count_282_pad;
  wire [11:0] count_35_shl;
  wire [19:0] count_35_pad;
  wire [10:0] count_428_shl;
  wire [19:0] count_428_pad;
  wire [14:0] count_16_shl;
  wire [19:0] count_16_pad;
  wire [11:0] count_355_shl;
  wire [19:0] count_355_pad;
  wire  count_110_shl;
  wire [19:0] count_110_pad;
  wire [18:0] count_367_shl;
  wire [19:0] count_367_pad;
  wire [17:0] count_427_shl;
  wire [19:0] count_427_pad;
  wire [2:0] count_46_shl;
  wire [19:0] count_46_pad;
  wire [3:0] count_272_shl;
  wire [19:0] count_272_pad;
  wire [17:0] count_5_shl;
  wire [19:0] count_5_pad;
  wire [6:0] count_173_shl;
  wire [19:0] count_173_pad;
  wire [18:0] count_211_shl;
  wire [19:0] count_211_pad;
  wire [1:0] count_230_shl;
  wire [19:0] count_230_pad;
  wire [7:0] count_454_shl;
  wire [19:0] count_454_pad;
  wire [10:0] count_458_shl;
  wire [19:0] count_458_pad;
  wire [5:0] count_23_shl;
  wire [19:0] count_23_pad;
  wire [12:0] count_350_shl;
  wire [19:0] count_350_pad;
  wire [7:0] count_368_shl;
  wire [19:0] count_368_pad;
  wire [7:0] count_456_shl;
  wire [19:0] count_456_pad;
  wire [6:0] count_464_shl;
  wire [19:0] count_464_pad;
  wire [3:0] count_56_shl;
  wire [19:0] count_56_pad;
  wire [6:0] count_158_shl;
  wire [19:0] count_158_pad;
  wire [13:0] count_1_shl;
  wire [19:0] count_1_pad;
  wire [7:0] count_62_shl;
  wire [19:0] count_62_pad;
  wire [4:0] count_295_shl;
  wire [19:0] count_295_pad;
  wire [7:0] count_285_shl;
  wire [19:0] count_285_pad;
  wire [9:0] count_44_shl;
  wire [19:0] count_44_pad;
  wire [17:0] count_25_shl;
  wire [19:0] count_25_pad;
  wire [1:0] count_256_shl;
  wire [19:0] count_256_pad;
  wire [17:0] count_366_shl;
  wire [19:0] count_366_pad;
  wire [13:0] count_473_shl;
  wire [19:0] count_473_pad;
  wire [2:0] count_465_shl;
  wire [19:0] count_465_pad;
  wire [10:0] count_268_shl;
  wire [19:0] count_268_pad;
  wire [19:0] count_142_shl;
  wire [19:0] count_142_pad;
  wire [4:0] count_75_shl;
  wire [19:0] count_75_pad;
  wire [9:0] count_240_shl;
  wire [19:0] count_240_pad;
  wire [2:0] count_481_shl;
  wire [19:0] count_481_pad;
  wire [1:0] count_189_shl;
  wire [19:0] count_189_pad;
  wire [4:0] count_382_shl;
  wire [19:0] count_382_pad;
  wire [1:0] count_219_shl;
  wire [19:0] count_219_pad;
  wire  count_365_shl;
  wire [19:0] count_365_pad;
  wire [9:0] count_300_shl;
  wire [19:0] count_300_pad;
  wire [13:0] count_53_shl;
  wire [19:0] count_53_pad;
  wire [16:0] count_490_shl;
  wire [19:0] count_490_pad;
  wire [19:0] count_190_shl;
  wire [19:0] count_190_pad;
  wire [9:0] count_332_shl;
  wire [19:0] count_332_pad;
  wire [4:0] count_258_shl;
  wire [19:0] count_258_pad;
  wire [18:0] count_356_shl;
  wire [19:0] count_356_pad;
  wire [7:0] count_410_shl;
  wire [19:0] count_410_pad;
  wire [5:0] count_68_shl;
  wire [19:0] count_68_pad;
  wire [9:0] count_444_shl;
  wire [19:0] count_444_pad;
  wire [14:0] count_446_shl;
  wire [19:0] count_446_pad;
  wire [11:0] count_493_shl;
  wire [19:0] count_493_pad;
  wire [5:0] count_404_shl;
  wire [19:0] count_404_pad;
  wire [15:0] count_40_shl;
  wire [19:0] count_40_pad;
  wire [14:0] count_495_shl;
  wire [19:0] count_495_pad;
  wire [16:0] count_325_shl;
  wire [19:0] count_325_pad;
  wire  count_58_shl;
  wire [19:0] count_58_pad;
  wire [19:0] count_201_shl;
  wire [19:0] count_201_pad;
  wire [18:0] count_107_shl;
  wire [19:0] count_107_pad;
  wire [6:0] count_292_shl;
  wire [19:0] count_292_pad;
  wire [4:0] count_462_shl;
  wire [19:0] count_462_pad;
  wire  count_380_shl;
  wire [19:0] count_380_pad;
  wire [16:0] count_57_shl;
  wire [19:0] count_57_pad;
  wire [6:0] count_395_shl;
  wire [19:0] count_395_pad;
  wire [18:0] count_20_shl;
  wire [19:0] count_20_pad;
  wire [10:0] count_99_shl;
  wire [19:0] count_99_pad;
  wire [19:0] count_327_shl;
  wire [19:0] count_327_pad;
  wire [1:0] count_30_shl;
  wire [19:0] count_30_pad;
  wire [7:0] count_302_shl;
  wire [19:0] count_302_pad;
  wire [14:0] count_77_shl;
  wire [19:0] count_77_pad;
  wire [6:0] count_439_shl;
  wire [19:0] count_439_pad;
  wire  count_409_shl;
  wire [19:0] count_409_pad;
  wire [8:0] count_443_shl;
  wire [19:0] count_443_pad;
  wire [10:0] count_143_shl;
  wire [19:0] count_143_pad;
  wire [5:0] count_165_shl;
  wire [19:0] count_165_pad;
  wire [17:0] count_81_shl;
  wire [19:0] count_81_pad;
  wire [19:0] count_346_shl;
  wire [19:0] count_346_pad;
  wire [6:0] count_314_shl;
  wire [19:0] count_314_pad;
  wire [5:0] count_196_shl;
  wire [19:0] count_196_pad;
  wire [2:0] count_262_shl;
  wire [19:0] count_262_pad;
  wire [14:0] count_402_shl;
  wire [19:0] count_402_pad;
  wire [18:0] count_87_shl;
  wire [19:0] count_87_pad;
  wire [5:0] count_29_shl;
  wire [19:0] count_29_pad;
  wire [13:0] count_126_shl;
  wire [19:0] count_126_pad;
  wire [6:0] count_318_shl;
  wire [19:0] count_318_pad;
  wire [2:0] count_66_shl;
  wire [19:0] count_66_pad;
  wire [1:0] count_163_shl;
  wire [19:0] count_163_pad;
  wire [4:0] count_175_shl;
  wire [19:0] count_175_pad;
  wire [14:0] count_71_shl;
  wire [19:0] count_71_pad;
  wire [9:0] count_80_shl;
  wire [19:0] count_80_pad;
  wire  count_252_shl;
  wire [19:0] count_252_pad;
  wire [6:0] count_28_shl;
  wire [19:0] count_28_pad;
  wire [17:0] count_502_shl;
  wire [19:0] count_502_pad;
  wire [19:0] count_459_shl;
  wire [19:0] count_459_pad;
  wire [15:0] count_141_shl;
  wire [19:0] count_141_pad;
  wire [16:0] count_405_shl;
  wire [19:0] count_405_pad;
  wire [3:0] count_511_shl;
  wire [19:0] count_511_pad;
  wire [7:0] count_254_shl;
  wire [19:0] count_254_pad;
  wire [15:0] count_476_shl;
  wire [19:0] count_476_pad;
  wire [2:0] count_97_shl;
  wire [19:0] count_97_pad;
  wire [3:0] count_448_shl;
  wire [19:0] count_448_pad;
  wire [12:0] count_193_shl;
  wire [19:0] count_193_pad;
  wire [16:0] count_260_shl;
  wire [19:0] count_260_pad;
  wire [18:0] count_303_shl;
  wire [19:0] count_303_pad;
  wire [6:0] count_177_shl;
  wire [19:0] count_177_pad;
  wire [6:0] count_470_shl;
  wire [19:0] count_470_pad;
  wire [8:0] count_146_shl;
  wire [19:0] count_146_pad;
  wire  count_309_shl;
  wire [19:0] count_309_pad;
  wire [12:0] count_213_shl;
  wire [19:0] count_213_pad;
  wire [17:0] count_343_shl;
  wire [19:0] count_343_pad;
  wire [16:0] count_468_shl;
  wire [19:0] count_468_pad;
  wire [7:0] count_429_shl;
  wire [19:0] count_429_pad;
  wire [12:0] count_244_shl;
  wire [19:0] count_244_pad;
  wire [19:0] count_69_shl;
  wire [19:0] count_69_pad;
  wire [19:0] count_460_shl;
  wire [19:0] count_460_pad;
  wire  count_370_shl;
  wire [19:0] count_370_pad;
  wire [10:0] count_125_shl;
  wire [19:0] count_125_pad;
  wire [12:0] count_290_shl;
  wire [19:0] count_290_pad;
  wire  count_128_shl;
  wire [19:0] count_128_pad;
  wire [13:0] count_407_shl;
  wire [19:0] count_407_pad;
  wire [9:0] count_198_shl;
  wire [19:0] count_198_pad;
  wire [4:0] count_140_shl;
  wire [19:0] count_140_pad;
  wire [9:0] count_512_shl;
  wire [19:0] count_512_pad;
  wire [9:0] count_440_shl;
  wire [19:0] count_440_pad;
  wire [4:0] count_362_shl;
  wire [19:0] count_362_pad;
  wire [12:0] count_480_shl;
  wire [19:0] count_480_pad;
  wire [10:0] count_109_shl;
  wire [19:0] count_109_pad;
  wire [10:0] count_171_shl;
  wire [19:0] count_171_pad;
  wire [18:0] count_414_shl;
  wire [19:0] count_414_pad;
  wire [17:0] count_267_shl;
  wire [19:0] count_267_pad;
  wire [13:0] count_484_shl;
  wire [19:0] count_484_pad;
  wire [8:0] count_278_shl;
  wire [19:0] count_278_pad;
  wire [9:0] count_39_shl;
  wire [19:0] count_39_pad;
  wire [9:0] count_360_shl;
  wire [19:0] count_360_pad;
  wire [1:0] count_14_shl;
  wire [19:0] count_14_pad;
  wire [10:0] count_336_shl;
  wire [19:0] count_336_pad;
  wire [8:0] count_108_shl;
  wire [19:0] count_108_pad;
  wire [8:0] count_45_shl;
  wire [19:0] count_45_pad;
  wire [5:0] count_275_shl;
  wire [19:0] count_275_pad;
  wire [7:0] count_413_shl;
  wire [19:0] count_413_pad;
  wire [9:0] count_52_shl;
  wire [19:0] count_52_pad;
  wire [9:0] count_41_shl;
  wire [19:0] count_41_pad;
  wire [13:0] count_328_shl;
  wire [19:0] count_328_pad;
  wire [16:0] count_82_shl;
  wire [19:0] count_82_pad;
  wire [18:0] count_4_shl;
  wire [19:0] count_4_pad;
  wire [19:0] count_299_shl;
  wire [19:0] count_299_pad;
  wire [1:0] count_286_shl;
  wire [19:0] count_286_pad;
  wire [1:0] count_510_shl;
  wire [19:0] count_510_pad;
  wire [11:0] count_96_shl;
  wire [19:0] count_96_pad;
  wire [7:0] count_203_shl;
  wire [19:0] count_203_pad;
  wire [15:0] count_452_shl;
  wire [19:0] count_452_pad;
  wire [13:0] count_150_shl;
  wire [19:0] count_150_pad;
  wire [2:0] count_385_shl;
  wire [19:0] count_385_pad;
  wire [7:0] count_156_shl;
  wire [19:0] count_156_pad;
  wire [15:0] count_169_shl;
  wire [19:0] count_169_pad;
  wire [10:0] count_132_shl;
  wire [19:0] count_132_pad;
  wire [12:0] count_225_shl;
  wire [19:0] count_225_pad;
  wire [19:0] count_341_shl;
  wire [19:0] count_341_pad;
  wire [2:0] count_377_shl;
  wire [19:0] count_377_pad;
  wire [6:0] count_114_shl;
  wire [19:0] count_114_pad;
  wire [7:0] count_294_shl;
  wire [19:0] count_294_pad;
  wire [12:0] count_79_shl;
  wire [19:0] count_79_pad;
  wire [15:0] count_60_shl;
  wire [19:0] count_60_pad;
  wire [1:0] count_86_shl;
  wire [19:0] count_86_pad;
  wire [14:0] count_399_shl;
  wire [19:0] count_399_pad;
  wire [15:0] count_279_shl;
  wire [19:0] count_279_pad;
  wire [15:0] count_239_shl;
  wire [19:0] count_239_pad;
  wire [12:0] count_13_shl;
  wire [19:0] count_13_pad;
  wire [16:0] count_337_shl;
  wire [19:0] count_337_pad;
  wire [5:0] count_19_shl;
  wire [19:0] count_19_pad;
  wire [9:0] count_334_shl;
  wire [19:0] count_334_pad;
  wire [16:0] count_17_shl;
  wire [19:0] count_17_pad;
  wire [5:0] count_72_shl;
  wire [19:0] count_72_pad;
  wire [14:0] count_94_shl;
  wire [19:0] count_94_pad;
  wire [5:0] count_419_shl;
  wire [19:0] count_419_pad;
  wire  count_176_shl;
  wire [19:0] count_176_pad;
  wire [11:0] count_210_shl;
  wire [19:0] count_210_pad;
  wire [14:0] count_78_shl;
  wire [19:0] count_78_pad;
  wire [17:0] count_104_shl;
  wire [19:0] count_104_pad;
  wire [19:0] count_507_shl;
  wire [19:0] count_507_pad;
  wire [17:0] count_287_shl;
  wire [19:0] count_287_pad;
  wire  count_208_shl;
  wire [19:0] count_208_pad;
  wire [9:0] count_345_shl;
  wire [19:0] count_345_pad;
  wire [14:0] count_311_shl;
  wire [19:0] count_311_pad;
  wire [3:0] count_178_shl;
  wire [19:0] count_178_pad;
  wire [6:0] count_89_shl;
  wire [19:0] count_89_pad;
  wire [17:0] count_266_shl;
  wire [19:0] count_266_pad;
  wire [2:0] count_238_shl;
  wire [19:0] count_238_pad;
  wire [5:0] count_206_shl;
  wire [19:0] count_206_pad;
  wire [18:0] count_103_shl;
  wire [19:0] count_103_pad;
  wire [15:0] count_85_shl;
  wire [19:0] count_85_pad;
  wire [15:0] count_138_shl;
  wire [19:0] count_138_pad;
  wire [18:0] count_392_shl;
  wire [19:0] count_392_pad;
  wire [16:0] count_271_shl;
  wire [19:0] count_271_pad;
  wire [15:0] count_445_shl;
  wire [19:0] count_445_pad;
  wire [10:0] count_431_shl;
  wire [19:0] count_431_pad;
  wire [14:0] count_220_shl;
  wire [19:0] count_220_pad;
  wire [9:0] count_160_shl;
  wire [19:0] count_160_pad;
  wire [11:0] count_183_shl;
  wire [19:0] count_183_pad;
  wire [13:0] count_436_shl;
  wire [19:0] count_436_pad;
  wire [19:0] count_226_shl;
  wire [19:0] count_226_pad;
  wire [16:0] count_136_shl;
  wire [19:0] count_136_pad;
  wire [18:0] count_42_shl;
  wire [19:0] count_42_pad;
  wire  count_351_shl;
  wire [19:0] count_351_pad;
  wire [17:0] count_261_shl;
  wire [19:0] count_261_pad;
  wire [4:0] count_221_shl;
  wire [19:0] count_221_pad;
  wire  count_152_shl;
  wire [19:0] count_152_pad;
  wire [7:0] count_505_shl;
  wire [19:0] count_505_pad;
  wire [9:0] count_36_shl;
  wire [19:0] count_36_pad;
  wire [13:0] count_232_shl;
  wire [19:0] count_232_pad;
  wire [5:0] count_479_shl;
  wire [19:0] count_479_pad;
  wire [19:0] count_34_shl;
  wire [19:0] count_34_pad;
  wire [4:0] count_291_shl;
  wire [19:0] count_291_pad;
  wire [11:0] count_246_shl;
  wire [19:0] count_246_pad;
  wire [15:0] count_9_shl;
  wire [19:0] count_9_pad;
  wire [3:0] count_98_shl;
  wire [19:0] count_98_pad;
  wire [1:0] count_364_shl;
  wire [19:0] count_364_pad;
  wire [14:0] count_451_shl;
  wire [19:0] count_451_pad;
  wire [16:0] count_426_shl;
  wire [19:0] count_426_pad;
  wire [1:0] count_492_shl;
  wire [19:0] count_492_pad;
  wire [4:0] count_281_shl;
  wire [19:0] count_281_pad;
  wire  count_494_shl;
  wire [19:0] count_494_pad;
  wire [13:0] count_340_shl;
  wire [19:0] count_340_pad;
  wire [9:0] count_179_shl;
  wire [19:0] count_179_pad;
  wire [16:0] count_250_shl;
  wire [19:0] count_250_pad;
  wire [10:0] count_249_shl;
  wire [19:0] count_249_pad;
  wire [8:0] count_59_shl;
  wire [19:0] count_59_pad;
  wire [6:0] count_320_shl;
  wire [19:0] count_320_pad;
  wire [16:0] count_321_shl;
  wire [19:0] count_321_pad;
  wire [14:0] count_449_shl;
  wire [19:0] count_449_pad;
  wire [8:0] count_2_shl;
  wire [19:0] count_2_pad;
  wire [11:0] count_496_shl;
  wire [19:0] count_496_pad;
  wire [2:0] count_188_shl;
  wire [19:0] count_188_pad;
  wire [13:0] count_466_shl;
  wire [19:0] count_466_pad;
  wire [18:0] count_212_shl;
  wire [19:0] count_212_pad;
  wire [18:0] count_11_shl;
  wire [19:0] count_11_pad;
  wire [16:0] count_55_shl;
  wire [19:0] count_55_pad;
  wire [2:0] count_119_shl;
  wire [19:0] count_119_pad;
  wire [10:0] count_149_shl;
  wire [19:0] count_149_pad;
  wire [9:0] count_450_shl;
  wire [19:0] count_450_pad;
  wire [11:0] count_32_shl;
  wire [19:0] count_32_pad;
  wire [19:0] count_319_shl;
  wire [19:0] count_319_pad;
  wire [1:0] count_384_shl;
  wire [19:0] count_384_pad;
  wire [9:0] count_162_shl;
  wire [19:0] count_162_pad;
  wire [14:0] count_231_shl;
  wire [19:0] count_231_pad;
  wire [8:0] count_63_shl;
  wire [19:0] count_63_pad;
  wire [5:0] count_489_shl;
  wire [19:0] count_489_pad;
  wire [4:0] count_509_shl;
  wire [19:0] count_509_pad;
  wire [1:0] count_133_shl;
  wire [19:0] count_133_pad;
  wire [10:0] count_415_shl;
  wire [19:0] count_415_pad;
  wire [7:0] count_323_shl;
  wire [19:0] count_323_pad;
  wire [2:0] count_289_shl;
  wire [19:0] count_289_pad;
  wire [1:0] count_342_shl;
  wire [19:0] count_342_pad;
  wire [5:0] count_408_shl;
  wire [19:0] count_408_pad;
  wire [8:0] count_22_shl;
  wire [19:0] count_22_pad;
  wire [9:0] count_308_shl;
  wire [19:0] count_308_pad;
  wire [15:0] count_424_shl;
  wire [19:0] count_424_pad;
  wire [2:0] count_353_shl;
  wire [19:0] count_353_pad;
  wire [3:0] count_217_shl;
  wire [19:0] count_217_pad;
  wire [2:0] count_497_shl;
  wire [19:0] count_497_pad;
  wire [12:0] count_430_shl;
  wire [19:0] count_430_pad;
  wire [4:0] count_369_shl;
  wire [19:0] count_369_pad;
  wire [12:0] count_463_shl;
  wire [19:0] count_463_pad;
  wire  count_389_shl;
  wire [19:0] count_389_pad;
  wire [3:0] count_499_shl;
  wire [19:0] count_499_pad;
  wire [13:0] count_315_shl;
  wire [19:0] count_315_pad;
  wire [5:0] count_113_shl;
  wire [19:0] count_113_pad;
  wire [12:0] count_506_shl;
  wire [19:0] count_506_pad;
  wire [19:0] count_257_shl;
  wire [19:0] count_257_pad;
  wire [10:0] count_12_shl;
  wire [19:0] count_12_pad;
  wire [18:0] count_397_shl;
  wire [19:0] count_397_pad;
  wire [10:0] count_326_shl;
  wire [19:0] count_326_pad;
  wire [13:0] count_469_shl;
  wire [19:0] count_469_pad;
  wire [17:0] count_316_shl;
  wire [19:0] count_316_pad;
  wire [11:0] count_248_shl;
  wire [19:0] count_248_pad;
  wire [12:0] r_first_shl;
  wire [19:0] r_first_pad;
  wire [18:0] count_390_shl;
  wire [19:0] count_390_pad;
  wire [19:0] count_277_shl;
  wire [19:0] count_277_pad;
  wire [7:0] count_269_shl;
  wire [19:0] count_269_pad;
  wire [10:0] count_218_shl;
  wire [19:0] count_218_pad;
  wire [13:0] count_115_shl;
  wire [19:0] count_115_pad;
  wire [14:0] count_166_shl;
  wire [19:0] count_166_pad;
  wire [18:0] count_487_shl;
  wire [19:0] count_487_pad;
  wire [2:0] count_192_shl;
  wire [19:0] count_192_pad;
  wire [19:0] count_508_shl;
  wire [19:0] count_508_pad;
  wire [8:0] count_358_shl;
  wire [19:0] count_358_pad;
  wire [15:0] count_416_shl;
  wire [19:0] count_416_pad;
  wire [9:0] count_151_shl;
  wire [19:0] count_151_pad;
  wire [12:0] count_354_shl;
  wire [19:0] count_354_pad;
  wire [19:0] count_21_shl;
  wire [19:0] count_21_pad;
  wire [18:0] r_holds_d_shl;
  wire [19:0] r_holds_d_pad;
  wire [18:0] count_339_shl;
  wire [19:0] count_339_pad;
  wire [15:0] count_111_shl;
  wire [19:0] count_111_pad;
  wire [17:0] count_18_shl;
  wire [19:0] count_18_pad;
  wire [17:0] count_425_shl;
  wire [19:0] count_425_pad;
  wire [19:0] count_455_shl;
  wire [19:0] count_455_pad;
  wire [4:0] count_437_shl;
  wire [19:0] count_437_pad;
  wire [16:0] count_245_shl;
  wire [19:0] count_245_pad;
  wire [10:0] count_116_shl;
  wire [19:0] count_116_pad;
  wire [3:0] count_194_shl;
  wire [19:0] count_194_pad;
  wire [5:0] count_127_shl;
  wire [19:0] count_127_pad;
  wire [6:0] count_137_shl;
  wire [19:0] count_137_pad;
  wire [2:0] count_483_shl;
  wire [19:0] count_483_pad;
  wire [3:0] count_159_shl;
  wire [19:0] count_159_pad;
  wire [15:0] count_301_shl;
  wire [19:0] count_301_pad;
  wire [18:0] count_215_shl;
  wire [19:0] count_215_pad;
  wire [9:0] count_288_shl;
  wire [19:0] count_288_pad;
  wire [5:0] count_54_shl;
  wire [19:0] count_54_pad;
  wire [18:0] count_27_shl;
  wire [19:0] count_27_pad;
  wire [16:0] count_161_shl;
  wire [19:0] count_161_pad;
  wire [1:0] count_106_shl;
  wire [19:0] count_106_pad;
  wire [7:0] count_485_shl;
  wire [19:0] count_485_pad;
  wire [3:0] count_259_shl;
  wire [19:0] count_259_pad;
  wire [11:0] count_264_shl;
  wire [19:0] count_264_pad;
  wire [9:0] count_91_shl;
  wire [19:0] count_91_pad;
  wire [1:0] count_84_shl;
  wire [19:0] count_84_pad;
  wire [3:0] count_312_shl;
  wire [19:0] count_312_pad;
  wire [3:0] count_207_shl;
  wire [19:0] count_207_pad;
  wire [7:0] count_172_shl;
  wire [19:0] count_172_pad;
  wire [11:0] count_253_shl;
  wire [19:0] count_253_pad;
  wire [12:0] count_148_shl;
  wire [19:0] count_148_pad;
  wire [1:0] count_228_shl;
  wire [19:0] count_228_pad;
  wire [3:0] count_10_shl;
  wire [19:0] count_10_pad;
  wire [9:0] count_322_shl;
  wire [19:0] count_322_pad;
  wire [9:0] count_363_shl;
  wire [19:0] count_363_pad;
  wire [11:0] count_48_shl;
  wire [19:0] count_48_pad;
  wire [16:0] count_236_shl;
  wire [19:0] count_236_pad;
  wire [16:0] count_205_shl;
  wire [19:0] count_205_pad;
  wire [15:0] count_191_shl;
  wire [19:0] count_191_pad;
  wire [4:0] count_338_shl;
  wire [19:0] count_338_pad;
  wire [16:0] count_276_shl;
  wire [19:0] count_276_pad;
  wire [2:0] count_475_shl;
  wire [19:0] count_475_pad;
  wire [15:0] count_24_shl;
  wire [19:0] count_24_pad;
  wire [16:0] count_387_shl;
  wire [19:0] count_387_pad;
  wire [8:0] count_438_shl;
  wire [19:0] count_438_pad;
  wire [3:0] count_472_shl;
  wire [19:0] count_472_pad;
  wire  count_167_shl;
  wire [19:0] count_167_pad;
  wire [2:0] count_233_shl;
  wire [19:0] count_233_pad;
  wire [6:0] count_185_shl;
  wire [19:0] count_185_pad;
  wire [12:0] count_135_shl;
  wire [19:0] count_135_pad;
  wire [18:0] count_197_shl;
  wire [19:0] count_197_pad;
  wire [19:0] count_273_shl;
  wire [19:0] count_273_pad;
  wire [14:0] count_441_shl;
  wire [19:0] count_441_pad;
  wire [1:0] count_88_shl;
  wire [19:0] count_88_pad;
  wire [13:0] count_471_shl;
  wire [19:0] count_471_pad;
  wire [9:0] count_147_shl;
  wire [19:0] count_147_pad;
  wire [17:0] count_412_shl;
  wire [19:0] count_412_pad;
  wire [18:0] count_488_shl;
  wire [19:0] count_488_pad;
  wire [8:0] count_486_shl;
  wire [19:0] count_486_pad;
  wire  count_298_shl;
  wire [19:0] count_298_pad;
  wire [8:0] count_442_shl;
  wire [19:0] count_442_pad;
  wire [9:0] count_73_shl;
  wire [19:0] count_73_pad;
  wire [13:0] count_237_shl;
  wire [19:0] count_237_pad;
  wire [12:0] count_435_shl;
  wire [19:0] count_435_pad;
  wire [6:0] count_6_shl;
  wire [19:0] count_6_pad;
  wire  count_361_shl;
  wire [19:0] count_361_pad;
  wire [1:0] count_15_shl;
  wire [19:0] count_15_pad;
  wire [12:0] count_388_shl;
  wire [19:0] count_388_pad;
  wire  count_164_shl;
  wire [19:0] count_164_pad;
  wire [3:0] count_255_shl;
  wire [19:0] count_255_pad;
  wire [18:0] count_306_shl;
  wire [19:0] count_306_pad;
  wire [19:0] count_381_shl;
  wire [19:0] count_381_pad;
  wire [6:0] count_130_shl;
  wire [19:0] count_130_pad;
  wire [18:0] count_145_shl;
  wire [19:0] count_145_pad;
  wire [5:0] count_8_shl;
  wire [19:0] count_8_pad;
  wire [6:0] count_224_shl;
  wire [19:0] count_224_pad;
  wire [12:0] count_349_shl;
  wire [19:0] count_349_pad;
  wire [18:0] count_375_shl;
  wire [19:0] count_375_pad;
  wire [18:0] count_457_shl;
  wire [19:0] count_457_pad;
  wire [8:0] b_delay_shl;
  wire [19:0] b_delay_pad;
  wire [15:0] count_181_shl;
  wire [19:0] count_181_pad;
  wire [13:0] count_170_shl;
  wire [19:0] count_170_pad;
  wire [7:0] count_3_shl;
  wire [19:0] count_3_pad;
  wire  count_461_shl;
  wire [19:0] count_461_pad;
  wire [11:0] count_102_shl;
  wire [19:0] count_102_pad;
  wire [2:0] count_134_shl;
  wire [19:0] count_134_pad;
  wire [17:0] count_234_shl;
  wire [19:0] count_234_pad;
  wire [19:0] count_335_shl;
  wire [19:0] count_335_pad;
  wire [12:0] count_95_shl;
  wire [19:0] count_95_pad;
  wire [6:0] count_374_shl;
  wire [19:0] count_374_pad;
  wire [2:0] count_49_shl;
  wire [19:0] count_49_pad;
  wire [8:0] count_100_shl;
  wire [19:0] count_100_pad;
  wire [6:0] count_283_shl;
  wire [19:0] count_283_pad;
  wire [17:0] count_90_shl;
  wire [19:0] count_90_pad;
  wire [9:0] count_155_shl;
  wire [19:0] count_155_pad;
  wire [1:0] count_274_shl;
  wire [19:0] count_274_pad;
  wire [13:0] count_83_shl;
  wire [19:0] count_83_pad;
  wire [11:0] count_112_shl;
  wire [19:0] count_112_pad;
  wire [12:0] count_433_shl;
  wire [19:0] count_433_pad;
  wire [1:0] count_93_shl;
  wire [19:0] count_93_pad;
  wire [3:0] count_65_shl;
  wire [19:0] count_65_pad;
  wire  count_235_shl;
  wire [19:0] count_235_pad;
  wire [3:0] count_371_shl;
  wire [19:0] count_371_pad;
  wire [5:0] count_122_shl;
  wire [19:0] count_122_pad;
  wire [13:0] count_247_shl;
  wire [19:0] count_247_pad;
  wire [11:0] count_157_shl;
  wire [19:0] count_157_pad;
  wire [6:0] count_180_shl;
  wire [19:0] count_180_pad;
  wire [13:0] count_347_shl;
  wire [19:0] count_347_pad;
  wire [16:0] count_251_shl;
  wire [19:0] count_251_pad;
  wire [15:0] count_200_shl;
  wire [19:0] count_200_pad;
  wire [8:0] count_187_shl;
  wire [19:0] count_187_pad;
  wire [5:0] count_432_shl;
  wire [19:0] count_432_pad;
  wire [2:0] count_123_shl;
  wire [19:0] count_123_pad;
  wire [3:0] count_418_shl;
  wire [19:0] count_418_pad;
  wire [4:0] count_406_shl;
  wire [19:0] count_406_pad;
  wire [18:0] count_241_shl;
  wire [19:0] count_241_pad;
  wire  count_33_shl;
  wire [19:0] count_33_pad;
  wire [12:0] count_324_shl;
  wire [19:0] count_324_pad;
  wire [5:0] count_105_shl;
  wire [19:0] count_105_pad;
  wire [1:0] count_92_shl;
  wire [19:0] count_92_pad;
  wire [5:0] count_7_shl;
  wire [19:0] count_7_pad;
  wire  count_214_shl;
  wire [19:0] count_214_pad;
  wire [11:0] count_379_shl;
  wire [19:0] count_379_pad;
  wire [7:0] count_359_shl;
  wire [19:0] count_359_pad;
  wire [16:0] doneAW_shl;
  wire [19:0] doneAW_pad;
  wire [6:0] count_144_shl;
  wire [19:0] count_144_pad;
  wire [18:0] count_396_shl;
  wire [19:0] count_396_pad;
  wire [4:0] count_376_shl;
  wire [19:0] count_376_pad;
  wire [18:0] count_504_shl;
  wire [19:0] count_504_pad;
  wire [6:0] count_124_shl;
  wire [19:0] count_124_pad;
  wire [13:0] count_500_shl;
  wire [19:0] count_500_pad;
  wire [18:0] count_209_shl;
  wire [19:0] count_209_pad;
  wire [19:0] count_348_shl;
  wire [19:0] count_348_pad;
  wire [16:0] count_344_shl;
  wire [19:0] count_344_pad;
  wire [16:0] count_76_shl;
  wire [19:0] count_76_pad;
  wire [5:0] count_265_shl;
  wire [19:0] count_265_pad;
  wire [7:0] count_453_shl;
  wire [19:0] count_453_pad;
  wire [9:0] count_47_shl;
  wire [19:0] count_47_pad;
  wire [2:0] count_43_shl;
  wire [19:0] count_43_pad;
  wire [5:0] count_74_shl;
  wire [19:0] count_74_pad;
  wire [6:0] count_491_shl;
  wire [19:0] count_491_pad;
  wire [9:0] count_478_shl;
  wire [19:0] count_478_pad;
  wire [6:0] count_243_shl;
  wire [19:0] count_243_pad;
  wire  count_174_shl;
  wire [19:0] count_174_pad;
  wire [19:0] TLToAXI4_xor255;
  wire [19:0] TLToAXI4_xor256;
  wire [19:0] TLToAXI4_xor127;
  wire [19:0] TLToAXI4_xor257;
  wire [19:0] TLToAXI4_xor258;
  wire [19:0] TLToAXI4_xor128;
  wire [19:0] TLToAXI4_xor63;
  wire [19:0] TLToAXI4_xor259;
  wire [19:0] TLToAXI4_xor260;
  wire [19:0] TLToAXI4_xor129;
  wire [19:0] TLToAXI4_xor261;
  wire [19:0] TLToAXI4_xor262;
  wire [19:0] TLToAXI4_xor130;
  wire [19:0] TLToAXI4_xor64;
  wire [19:0] TLToAXI4_xor31;
  wire [19:0] TLToAXI4_xor263;
  wire [19:0] TLToAXI4_xor264;
  wire [19:0] TLToAXI4_xor131;
  wire [19:0] TLToAXI4_xor265;
  wire [19:0] TLToAXI4_xor266;
  wire [19:0] TLToAXI4_xor132;
  wire [19:0] TLToAXI4_xor65;
  wire [19:0] TLToAXI4_xor267;
  wire [19:0] TLToAXI4_xor268;
  wire [19:0] TLToAXI4_xor133;
  wire [19:0] TLToAXI4_xor269;
  wire [19:0] TLToAXI4_xor270;
  wire [19:0] TLToAXI4_xor134;
  wire [19:0] TLToAXI4_xor66;
  wire [19:0] TLToAXI4_xor32;
  wire [19:0] TLToAXI4_xor15;
  wire [19:0] TLToAXI4_xor271;
  wire [19:0] TLToAXI4_xor272;
  wire [19:0] TLToAXI4_xor135;
  wire [19:0] TLToAXI4_xor273;
  wire [19:0] TLToAXI4_xor274;
  wire [19:0] TLToAXI4_xor136;
  wire [19:0] TLToAXI4_xor67;
  wire [19:0] TLToAXI4_xor275;
  wire [19:0] TLToAXI4_xor276;
  wire [19:0] TLToAXI4_xor137;
  wire [19:0] TLToAXI4_xor277;
  wire [19:0] TLToAXI4_xor278;
  wire [19:0] TLToAXI4_xor138;
  wire [19:0] TLToAXI4_xor68;
  wire [19:0] TLToAXI4_xor33;
  wire [19:0] TLToAXI4_xor279;
  wire [19:0] TLToAXI4_xor280;
  wire [19:0] TLToAXI4_xor139;
  wire [19:0] TLToAXI4_xor281;
  wire [19:0] TLToAXI4_xor282;
  wire [19:0] TLToAXI4_xor140;
  wire [19:0] TLToAXI4_xor69;
  wire [19:0] TLToAXI4_xor283;
  wire [19:0] TLToAXI4_xor284;
  wire [19:0] TLToAXI4_xor141;
  wire [19:0] TLToAXI4_xor285;
  wire [19:0] TLToAXI4_xor286;
  wire [19:0] TLToAXI4_xor142;
  wire [19:0] TLToAXI4_xor70;
  wire [19:0] TLToAXI4_xor34;
  wire [19:0] TLToAXI4_xor16;
  wire [19:0] TLToAXI4_xor7;
  wire [19:0] TLToAXI4_xor287;
  wire [19:0] TLToAXI4_xor288;
  wire [19:0] TLToAXI4_xor143;
  wire [19:0] TLToAXI4_xor289;
  wire [19:0] TLToAXI4_xor290;
  wire [19:0] TLToAXI4_xor144;
  wire [19:0] TLToAXI4_xor71;
  wire [19:0] TLToAXI4_xor291;
  wire [19:0] TLToAXI4_xor292;
  wire [19:0] TLToAXI4_xor145;
  wire [19:0] TLToAXI4_xor293;
  wire [19:0] TLToAXI4_xor294;
  wire [19:0] TLToAXI4_xor146;
  wire [19:0] TLToAXI4_xor72;
  wire [19:0] TLToAXI4_xor35;
  wire [19:0] TLToAXI4_xor295;
  wire [19:0] TLToAXI4_xor296;
  wire [19:0] TLToAXI4_xor147;
  wire [19:0] TLToAXI4_xor297;
  wire [19:0] TLToAXI4_xor298;
  wire [19:0] TLToAXI4_xor148;
  wire [19:0] TLToAXI4_xor73;
  wire [19:0] TLToAXI4_xor299;
  wire [19:0] TLToAXI4_xor300;
  wire [19:0] TLToAXI4_xor149;
  wire [19:0] TLToAXI4_xor301;
  wire [19:0] TLToAXI4_xor302;
  wire [19:0] TLToAXI4_xor150;
  wire [19:0] TLToAXI4_xor74;
  wire [19:0] TLToAXI4_xor36;
  wire [19:0] TLToAXI4_xor17;
  wire [19:0] TLToAXI4_xor303;
  wire [19:0] TLToAXI4_xor304;
  wire [19:0] TLToAXI4_xor151;
  wire [19:0] TLToAXI4_xor305;
  wire [19:0] TLToAXI4_xor306;
  wire [19:0] TLToAXI4_xor152;
  wire [19:0] TLToAXI4_xor75;
  wire [19:0] TLToAXI4_xor307;
  wire [19:0] TLToAXI4_xor308;
  wire [19:0] TLToAXI4_xor153;
  wire [19:0] TLToAXI4_xor309;
  wire [19:0] TLToAXI4_xor310;
  wire [19:0] TLToAXI4_xor154;
  wire [19:0] TLToAXI4_xor76;
  wire [19:0] TLToAXI4_xor37;
  wire [19:0] TLToAXI4_xor311;
  wire [19:0] TLToAXI4_xor312;
  wire [19:0] TLToAXI4_xor155;
  wire [19:0] TLToAXI4_xor313;
  wire [19:0] TLToAXI4_xor314;
  wire [19:0] TLToAXI4_xor156;
  wire [19:0] TLToAXI4_xor77;
  wire [19:0] TLToAXI4_xor315;
  wire [19:0] TLToAXI4_xor316;
  wire [19:0] TLToAXI4_xor157;
  wire [19:0] TLToAXI4_xor317;
  wire [19:0] TLToAXI4_xor638;
  wire [19:0] TLToAXI4_xor318;
  wire [19:0] TLToAXI4_xor158;
  wire [19:0] TLToAXI4_xor78;
  wire [19:0] TLToAXI4_xor38;
  wire [19:0] TLToAXI4_xor18;
  wire [19:0] TLToAXI4_xor8;
  wire [19:0] TLToAXI4_xor3;
  wire [19:0] TLToAXI4_xor319;
  wire [19:0] TLToAXI4_xor320;
  wire [19:0] TLToAXI4_xor159;
  wire [19:0] TLToAXI4_xor321;
  wire [19:0] TLToAXI4_xor322;
  wire [19:0] TLToAXI4_xor160;
  wire [19:0] TLToAXI4_xor79;
  wire [19:0] TLToAXI4_xor323;
  wire [19:0] TLToAXI4_xor324;
  wire [19:0] TLToAXI4_xor161;
  wire [19:0] TLToAXI4_xor325;
  wire [19:0] TLToAXI4_xor326;
  wire [19:0] TLToAXI4_xor162;
  wire [19:0] TLToAXI4_xor80;
  wire [19:0] TLToAXI4_xor39;
  wire [19:0] TLToAXI4_xor327;
  wire [19:0] TLToAXI4_xor328;
  wire [19:0] TLToAXI4_xor163;
  wire [19:0] TLToAXI4_xor329;
  wire [19:0] TLToAXI4_xor330;
  wire [19:0] TLToAXI4_xor164;
  wire [19:0] TLToAXI4_xor81;
  wire [19:0] TLToAXI4_xor331;
  wire [19:0] TLToAXI4_xor332;
  wire [19:0] TLToAXI4_xor165;
  wire [19:0] TLToAXI4_xor333;
  wire [19:0] TLToAXI4_xor334;
  wire [19:0] TLToAXI4_xor166;
  wire [19:0] TLToAXI4_xor82;
  wire [19:0] TLToAXI4_xor40;
  wire [19:0] TLToAXI4_xor19;
  wire [19:0] TLToAXI4_xor335;
  wire [19:0] TLToAXI4_xor336;
  wire [19:0] TLToAXI4_xor167;
  wire [19:0] TLToAXI4_xor337;
  wire [19:0] TLToAXI4_xor338;
  wire [19:0] TLToAXI4_xor168;
  wire [19:0] TLToAXI4_xor83;
  wire [19:0] TLToAXI4_xor339;
  wire [19:0] TLToAXI4_xor340;
  wire [19:0] TLToAXI4_xor169;
  wire [19:0] TLToAXI4_xor341;
  wire [19:0] TLToAXI4_xor342;
  wire [19:0] TLToAXI4_xor170;
  wire [19:0] TLToAXI4_xor84;
  wire [19:0] TLToAXI4_xor41;
  wire [19:0] TLToAXI4_xor343;
  wire [19:0] TLToAXI4_xor344;
  wire [19:0] TLToAXI4_xor171;
  wire [19:0] TLToAXI4_xor345;
  wire [19:0] TLToAXI4_xor346;
  wire [19:0] TLToAXI4_xor172;
  wire [19:0] TLToAXI4_xor85;
  wire [19:0] TLToAXI4_xor347;
  wire [19:0] TLToAXI4_xor348;
  wire [19:0] TLToAXI4_xor173;
  wire [19:0] TLToAXI4_xor349;
  wire [19:0] TLToAXI4_xor350;
  wire [19:0] TLToAXI4_xor174;
  wire [19:0] TLToAXI4_xor86;
  wire [19:0] TLToAXI4_xor42;
  wire [19:0] TLToAXI4_xor20;
  wire [19:0] TLToAXI4_xor9;
  wire [19:0] TLToAXI4_xor351;
  wire [19:0] TLToAXI4_xor352;
  wire [19:0] TLToAXI4_xor175;
  wire [19:0] TLToAXI4_xor353;
  wire [19:0] TLToAXI4_xor354;
  wire [19:0] TLToAXI4_xor176;
  wire [19:0] TLToAXI4_xor87;
  wire [19:0] TLToAXI4_xor355;
  wire [19:0] TLToAXI4_xor356;
  wire [19:0] TLToAXI4_xor177;
  wire [19:0] TLToAXI4_xor357;
  wire [19:0] TLToAXI4_xor358;
  wire [19:0] TLToAXI4_xor178;
  wire [19:0] TLToAXI4_xor88;
  wire [19:0] TLToAXI4_xor43;
  wire [19:0] TLToAXI4_xor359;
  wire [19:0] TLToAXI4_xor360;
  wire [19:0] TLToAXI4_xor179;
  wire [19:0] TLToAXI4_xor361;
  wire [19:0] TLToAXI4_xor362;
  wire [19:0] TLToAXI4_xor180;
  wire [19:0] TLToAXI4_xor89;
  wire [19:0] TLToAXI4_xor363;
  wire [19:0] TLToAXI4_xor364;
  wire [19:0] TLToAXI4_xor181;
  wire [19:0] TLToAXI4_xor365;
  wire [19:0] TLToAXI4_xor366;
  wire [19:0] TLToAXI4_xor182;
  wire [19:0] TLToAXI4_xor90;
  wire [19:0] TLToAXI4_xor44;
  wire [19:0] TLToAXI4_xor21;
  wire [19:0] TLToAXI4_xor367;
  wire [19:0] TLToAXI4_xor368;
  wire [19:0] TLToAXI4_xor183;
  wire [19:0] TLToAXI4_xor369;
  wire [19:0] TLToAXI4_xor370;
  wire [19:0] TLToAXI4_xor184;
  wire [19:0] TLToAXI4_xor91;
  wire [19:0] TLToAXI4_xor371;
  wire [19:0] TLToAXI4_xor372;
  wire [19:0] TLToAXI4_xor185;
  wire [19:0] TLToAXI4_xor373;
  wire [19:0] TLToAXI4_xor374;
  wire [19:0] TLToAXI4_xor186;
  wire [19:0] TLToAXI4_xor92;
  wire [19:0] TLToAXI4_xor45;
  wire [19:0] TLToAXI4_xor375;
  wire [19:0] TLToAXI4_xor376;
  wire [19:0] TLToAXI4_xor187;
  wire [19:0] TLToAXI4_xor377;
  wire [19:0] TLToAXI4_xor378;
  wire [19:0] TLToAXI4_xor188;
  wire [19:0] TLToAXI4_xor93;
  wire [19:0] TLToAXI4_xor379;
  wire [19:0] TLToAXI4_xor380;
  wire [19:0] TLToAXI4_xor189;
  wire [19:0] TLToAXI4_xor381;
  wire [19:0] TLToAXI4_xor766;
  wire [19:0] TLToAXI4_xor382;
  wire [19:0] TLToAXI4_xor190;
  wire [19:0] TLToAXI4_xor94;
  wire [19:0] TLToAXI4_xor46;
  wire [19:0] TLToAXI4_xor22;
  wire [19:0] TLToAXI4_xor10;
  wire [19:0] TLToAXI4_xor4;
  wire [19:0] TLToAXI4_xor1;
  wire [19:0] TLToAXI4_xor383;
  wire [19:0] TLToAXI4_xor384;
  wire [19:0] TLToAXI4_xor191;
  wire [19:0] TLToAXI4_xor385;
  wire [19:0] TLToAXI4_xor386;
  wire [19:0] TLToAXI4_xor192;
  wire [19:0] TLToAXI4_xor95;
  wire [19:0] TLToAXI4_xor387;
  wire [19:0] TLToAXI4_xor388;
  wire [19:0] TLToAXI4_xor193;
  wire [19:0] TLToAXI4_xor389;
  wire [19:0] TLToAXI4_xor390;
  wire [19:0] TLToAXI4_xor194;
  wire [19:0] TLToAXI4_xor96;
  wire [19:0] TLToAXI4_xor47;
  wire [19:0] TLToAXI4_xor391;
  wire [19:0] TLToAXI4_xor392;
  wire [19:0] TLToAXI4_xor195;
  wire [19:0] TLToAXI4_xor393;
  wire [19:0] TLToAXI4_xor394;
  wire [19:0] TLToAXI4_xor196;
  wire [19:0] TLToAXI4_xor97;
  wire [19:0] TLToAXI4_xor395;
  wire [19:0] TLToAXI4_xor396;
  wire [19:0] TLToAXI4_xor197;
  wire [19:0] TLToAXI4_xor397;
  wire [19:0] TLToAXI4_xor398;
  wire [19:0] TLToAXI4_xor198;
  wire [19:0] TLToAXI4_xor98;
  wire [19:0] TLToAXI4_xor48;
  wire [19:0] TLToAXI4_xor23;
  wire [19:0] TLToAXI4_xor399;
  wire [19:0] TLToAXI4_xor400;
  wire [19:0] TLToAXI4_xor199;
  wire [19:0] TLToAXI4_xor401;
  wire [19:0] TLToAXI4_xor402;
  wire [19:0] TLToAXI4_xor200;
  wire [19:0] TLToAXI4_xor99;
  wire [19:0] TLToAXI4_xor403;
  wire [19:0] TLToAXI4_xor404;
  wire [19:0] TLToAXI4_xor201;
  wire [19:0] TLToAXI4_xor405;
  wire [19:0] TLToAXI4_xor406;
  wire [19:0] TLToAXI4_xor202;
  wire [19:0] TLToAXI4_xor100;
  wire [19:0] TLToAXI4_xor49;
  wire [19:0] TLToAXI4_xor407;
  wire [19:0] TLToAXI4_xor408;
  wire [19:0] TLToAXI4_xor203;
  wire [19:0] TLToAXI4_xor409;
  wire [19:0] TLToAXI4_xor410;
  wire [19:0] TLToAXI4_xor204;
  wire [19:0] TLToAXI4_xor101;
  wire [19:0] TLToAXI4_xor411;
  wire [19:0] TLToAXI4_xor412;
  wire [19:0] TLToAXI4_xor205;
  wire [19:0] TLToAXI4_xor413;
  wire [19:0] TLToAXI4_xor414;
  wire [19:0] TLToAXI4_xor206;
  wire [19:0] TLToAXI4_xor102;
  wire [19:0] TLToAXI4_xor50;
  wire [19:0] TLToAXI4_xor24;
  wire [19:0] TLToAXI4_xor11;
  wire [19:0] TLToAXI4_xor415;
  wire [19:0] TLToAXI4_xor416;
  wire [19:0] TLToAXI4_xor207;
  wire [19:0] TLToAXI4_xor417;
  wire [19:0] TLToAXI4_xor418;
  wire [19:0] TLToAXI4_xor208;
  wire [19:0] TLToAXI4_xor103;
  wire [19:0] TLToAXI4_xor419;
  wire [19:0] TLToAXI4_xor420;
  wire [19:0] TLToAXI4_xor209;
  wire [19:0] TLToAXI4_xor421;
  wire [19:0] TLToAXI4_xor422;
  wire [19:0] TLToAXI4_xor210;
  wire [19:0] TLToAXI4_xor104;
  wire [19:0] TLToAXI4_xor51;
  wire [19:0] TLToAXI4_xor423;
  wire [19:0] TLToAXI4_xor424;
  wire [19:0] TLToAXI4_xor211;
  wire [19:0] TLToAXI4_xor425;
  wire [19:0] TLToAXI4_xor426;
  wire [19:0] TLToAXI4_xor212;
  wire [19:0] TLToAXI4_xor105;
  wire [19:0] TLToAXI4_xor427;
  wire [19:0] TLToAXI4_xor428;
  wire [19:0] TLToAXI4_xor213;
  wire [19:0] TLToAXI4_xor429;
  wire [19:0] TLToAXI4_xor430;
  wire [19:0] TLToAXI4_xor214;
  wire [19:0] TLToAXI4_xor106;
  wire [19:0] TLToAXI4_xor52;
  wire [19:0] TLToAXI4_xor25;
  wire [19:0] TLToAXI4_xor431;
  wire [19:0] TLToAXI4_xor432;
  wire [19:0] TLToAXI4_xor215;
  wire [19:0] TLToAXI4_xor433;
  wire [19:0] TLToAXI4_xor434;
  wire [19:0] TLToAXI4_xor216;
  wire [19:0] TLToAXI4_xor107;
  wire [19:0] TLToAXI4_xor435;
  wire [19:0] TLToAXI4_xor436;
  wire [19:0] TLToAXI4_xor217;
  wire [19:0] TLToAXI4_xor437;
  wire [19:0] TLToAXI4_xor438;
  wire [19:0] TLToAXI4_xor218;
  wire [19:0] TLToAXI4_xor108;
  wire [19:0] TLToAXI4_xor53;
  wire [19:0] TLToAXI4_xor439;
  wire [19:0] TLToAXI4_xor440;
  wire [19:0] TLToAXI4_xor219;
  wire [19:0] TLToAXI4_xor441;
  wire [19:0] TLToAXI4_xor442;
  wire [19:0] TLToAXI4_xor220;
  wire [19:0] TLToAXI4_xor109;
  wire [19:0] TLToAXI4_xor443;
  wire [19:0] TLToAXI4_xor444;
  wire [19:0] TLToAXI4_xor221;
  wire [19:0] TLToAXI4_xor445;
  wire [19:0] TLToAXI4_xor894;
  wire [19:0] TLToAXI4_xor446;
  wire [19:0] TLToAXI4_xor222;
  wire [19:0] TLToAXI4_xor110;
  wire [19:0] TLToAXI4_xor54;
  wire [19:0] TLToAXI4_xor26;
  wire [19:0] TLToAXI4_xor12;
  wire [19:0] TLToAXI4_xor5;
  wire [19:0] TLToAXI4_xor447;
  wire [19:0] TLToAXI4_xor448;
  wire [19:0] TLToAXI4_xor223;
  wire [19:0] TLToAXI4_xor449;
  wire [19:0] TLToAXI4_xor450;
  wire [19:0] TLToAXI4_xor224;
  wire [19:0] TLToAXI4_xor111;
  wire [19:0] TLToAXI4_xor451;
  wire [19:0] TLToAXI4_xor452;
  wire [19:0] TLToAXI4_xor225;
  wire [19:0] TLToAXI4_xor453;
  wire [19:0] TLToAXI4_xor454;
  wire [19:0] TLToAXI4_xor226;
  wire [19:0] TLToAXI4_xor112;
  wire [19:0] TLToAXI4_xor55;
  wire [19:0] TLToAXI4_xor455;
  wire [19:0] TLToAXI4_xor456;
  wire [19:0] TLToAXI4_xor227;
  wire [19:0] TLToAXI4_xor457;
  wire [19:0] TLToAXI4_xor458;
  wire [19:0] TLToAXI4_xor228;
  wire [19:0] TLToAXI4_xor113;
  wire [19:0] TLToAXI4_xor459;
  wire [19:0] TLToAXI4_xor460;
  wire [19:0] TLToAXI4_xor229;
  wire [19:0] TLToAXI4_xor461;
  wire [19:0] TLToAXI4_xor462;
  wire [19:0] TLToAXI4_xor230;
  wire [19:0] TLToAXI4_xor114;
  wire [19:0] TLToAXI4_xor56;
  wire [19:0] TLToAXI4_xor27;
  wire [19:0] TLToAXI4_xor463;
  wire [19:0] TLToAXI4_xor464;
  wire [19:0] TLToAXI4_xor231;
  wire [19:0] TLToAXI4_xor465;
  wire [19:0] TLToAXI4_xor466;
  wire [19:0] TLToAXI4_xor232;
  wire [19:0] TLToAXI4_xor115;
  wire [19:0] TLToAXI4_xor467;
  wire [19:0] TLToAXI4_xor468;
  wire [19:0] TLToAXI4_xor233;
  wire [19:0] TLToAXI4_xor469;
  wire [19:0] TLToAXI4_xor470;
  wire [19:0] TLToAXI4_xor234;
  wire [19:0] TLToAXI4_xor116;
  wire [19:0] TLToAXI4_xor57;
  wire [19:0] TLToAXI4_xor471;
  wire [19:0] TLToAXI4_xor472;
  wire [19:0] TLToAXI4_xor235;
  wire [19:0] TLToAXI4_xor473;
  wire [19:0] TLToAXI4_xor474;
  wire [19:0] TLToAXI4_xor236;
  wire [19:0] TLToAXI4_xor117;
  wire [19:0] TLToAXI4_xor475;
  wire [19:0] TLToAXI4_xor476;
  wire [19:0] TLToAXI4_xor237;
  wire [19:0] TLToAXI4_xor477;
  wire [19:0] TLToAXI4_xor478;
  wire [19:0] TLToAXI4_xor238;
  wire [19:0] TLToAXI4_xor118;
  wire [19:0] TLToAXI4_xor58;
  wire [19:0] TLToAXI4_xor28;
  wire [19:0] TLToAXI4_xor13;
  wire [19:0] TLToAXI4_xor479;
  wire [19:0] TLToAXI4_xor480;
  wire [19:0] TLToAXI4_xor239;
  wire [19:0] TLToAXI4_xor481;
  wire [19:0] TLToAXI4_xor482;
  wire [19:0] TLToAXI4_xor240;
  wire [19:0] TLToAXI4_xor119;
  wire [19:0] TLToAXI4_xor483;
  wire [19:0] TLToAXI4_xor484;
  wire [19:0] TLToAXI4_xor241;
  wire [19:0] TLToAXI4_xor485;
  wire [19:0] TLToAXI4_xor486;
  wire [19:0] TLToAXI4_xor242;
  wire [19:0] TLToAXI4_xor120;
  wire [19:0] TLToAXI4_xor59;
  wire [19:0] TLToAXI4_xor487;
  wire [19:0] TLToAXI4_xor488;
  wire [19:0] TLToAXI4_xor243;
  wire [19:0] TLToAXI4_xor489;
  wire [19:0] TLToAXI4_xor490;
  wire [19:0] TLToAXI4_xor244;
  wire [19:0] TLToAXI4_xor121;
  wire [19:0] TLToAXI4_xor491;
  wire [19:0] TLToAXI4_xor492;
  wire [19:0] TLToAXI4_xor245;
  wire [19:0] TLToAXI4_xor493;
  wire [19:0] TLToAXI4_xor494;
  wire [19:0] TLToAXI4_xor246;
  wire [19:0] TLToAXI4_xor122;
  wire [19:0] TLToAXI4_xor60;
  wire [19:0] TLToAXI4_xor29;
  wire [19:0] TLToAXI4_xor495;
  wire [19:0] TLToAXI4_xor496;
  wire [19:0] TLToAXI4_xor247;
  wire [19:0] TLToAXI4_xor497;
  wire [19:0] TLToAXI4_xor498;
  wire [19:0] TLToAXI4_xor248;
  wire [19:0] TLToAXI4_xor123;
  wire [19:0] TLToAXI4_xor499;
  wire [19:0] TLToAXI4_xor500;
  wire [19:0] TLToAXI4_xor249;
  wire [19:0] TLToAXI4_xor501;
  wire [19:0] TLToAXI4_xor502;
  wire [19:0] TLToAXI4_xor250;
  wire [19:0] TLToAXI4_xor124;
  wire [19:0] TLToAXI4_xor61;
  wire [19:0] TLToAXI4_xor503;
  wire [19:0] TLToAXI4_xor504;
  wire [19:0] TLToAXI4_xor251;
  wire [19:0] TLToAXI4_xor505;
  wire [19:0] TLToAXI4_xor506;
  wire [19:0] TLToAXI4_xor252;
  wire [19:0] TLToAXI4_xor125;
  wire [19:0] TLToAXI4_xor507;
  wire [19:0] TLToAXI4_xor508;
  wire [19:0] TLToAXI4_xor253;
  wire [19:0] TLToAXI4_xor509;
  wire [19:0] TLToAXI4_xor1022;
  wire [19:0] TLToAXI4_xor510;
  wire [19:0] TLToAXI4_xor254;
  wire [19:0] TLToAXI4_xor126;
  wire [19:0] TLToAXI4_xor62;
  wire [19:0] TLToAXI4_xor30;
  wire [19:0] TLToAXI4_xor14;
  wire [19:0] TLToAXI4_xor6;
  wire [19:0] TLToAXI4_xor2;
  wire [19:0] TLToAXI4_xor0;
  wire [29:0] deq_sum;
  wire [29:0] queue_arw_deq_sum;
  Queue_12 deq ( // @[Decoupled.scala 361:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_data(deq_io_enq_bits_data),
    .io_enq_bits_strb(deq_io_enq_bits_strb),
    .io_enq_bits_last(deq_io_enq_bits_last),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_data(deq_io_deq_bits_data),
    .io_deq_bits_strb(deq_io_deq_bits_strb),
    .io_deq_bits_last(deq_io_deq_bits_last),
    .io_covSum(deq_io_covSum),
    .metaReset(deq_metaReset)
  );
  Queue_19 queue_arw_deq ( // @[Decoupled.scala 361:21]
    .clock(queue_arw_deq_clock),
    .reset(queue_arw_deq_reset),
    .io_enq_ready(queue_arw_deq_io_enq_ready),
    .io_enq_valid(queue_arw_deq_io_enq_valid),
    .io_enq_bits_id(queue_arw_deq_io_enq_bits_id),
    .io_enq_bits_addr(queue_arw_deq_io_enq_bits_addr),
    .io_enq_bits_len(queue_arw_deq_io_enq_bits_len),
    .io_enq_bits_size(queue_arw_deq_io_enq_bits_size),
    .io_enq_bits_cache(queue_arw_deq_io_enq_bits_cache),
    .io_enq_bits_prot(queue_arw_deq_io_enq_bits_prot),
    .io_enq_bits_echo_tl_state_size(queue_arw_deq_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(queue_arw_deq_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_wen(queue_arw_deq_io_enq_bits_wen),
    .io_deq_ready(queue_arw_deq_io_deq_ready),
    .io_deq_valid(queue_arw_deq_io_deq_valid),
    .io_deq_bits_id(queue_arw_deq_io_deq_bits_id),
    .io_deq_bits_addr(queue_arw_deq_io_deq_bits_addr),
    .io_deq_bits_len(queue_arw_deq_io_deq_bits_len),
    .io_deq_bits_size(queue_arw_deq_io_deq_bits_size),
    .io_deq_bits_burst(queue_arw_deq_io_deq_bits_burst),
    .io_deq_bits_lock(queue_arw_deq_io_deq_bits_lock),
    .io_deq_bits_cache(queue_arw_deq_io_deq_bits_cache),
    .io_deq_bits_prot(queue_arw_deq_io_deq_bits_prot),
    .io_deq_bits_qos(queue_arw_deq_io_deq_bits_qos),
    .io_deq_bits_echo_tl_state_size(queue_arw_deq_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(queue_arw_deq_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_wen(queue_arw_deq_io_deq_bits_wen),
    .io_covSum(queue_arw_deq_io_covSum),
    .metaReset(queue_arw_deq_metaReset)
  );
  assign auto_in_a_ready = ~stall & _bundleIn_0_a_ready_T_3; // @[ToAXI4.scala 196:28]
  assign auto_in_d_valid = r_wins ? auto_out_r_valid : auto_out_b_valid; // @[ToAXI4.scala 219:24]
  assign auto_in_d_bits_opcode = r_wins ? 3'h1 : 3'h0; // @[ToAXI4.scala 237:23]
  assign auto_in_d_bits_size = r_wins ? r_d_size : b_d_size; // @[ToAXI4.scala 237:23]
  assign auto_in_d_bits_source = r_wins ? auto_out_r_bits_echo_tl_state_source : auto_out_b_bits_echo_tl_state_source; // @[ToAXI4.scala 237:23]
  assign auto_in_d_bits_denied = r_wins ? _GEN_1029 : b_denied; // @[ToAXI4.scala 237:23]
  assign auto_in_d_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = r_wins & r_d_corrupt; // @[ToAXI4.scala 237:23]
  assign auto_out_aw_valid = queue_arw_valid & queue_arw_bits_wen; // @[ToAXI4.scala 156:39]
  assign auto_out_aw_bits_id = queue_arw_deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_addr = queue_arw_deq_io_deq_bits_addr; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_len = queue_arw_deq_io_deq_bits_len; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_size = queue_arw_deq_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_burst = queue_arw_deq_io_deq_bits_burst; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_lock = queue_arw_deq_io_deq_bits_lock; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_cache = queue_arw_deq_io_deq_bits_cache; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_prot = queue_arw_deq_io_deq_bits_prot; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_qos = queue_arw_deq_io_deq_bits_qos; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_echo_tl_state_size = queue_arw_deq_io_deq_bits_echo_tl_state_size; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_echo_tl_state_source = queue_arw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_w_valid = deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  assign auto_out_w_bits_data = deq_io_deq_bits_data; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_w_bits_strb = deq_io_deq_bits_strb; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_w_bits_last = deq_io_deq_bits_last; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_b_ready = auto_in_d_ready & ~r_wins; // @[ToAXI4.scala 218:33]
  assign auto_out_ar_valid = queue_arw_valid & ~queue_arw_bits_wen; // @[ToAXI4.scala 155:39]
  assign auto_out_ar_bits_id = queue_arw_deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_addr = queue_arw_deq_io_deq_bits_addr; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_len = queue_arw_deq_io_deq_bits_len; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_size = queue_arw_deq_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_burst = queue_arw_deq_io_deq_bits_burst; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_lock = queue_arw_deq_io_deq_bits_lock; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_cache = queue_arw_deq_io_deq_bits_cache; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_prot = queue_arw_deq_io_deq_bits_prot; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_qos = queue_arw_deq_io_deq_bits_qos; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_echo_tl_state_size = queue_arw_deq_io_deq_bits_echo_tl_state_size; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_echo_tl_state_source = queue_arw_deq_io_deq_bits_echo_tl_state_source; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_r_ready = auto_in_d_ready & r_wins; // @[ToAXI4.scala 217:33]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = _out_arw_valid_T_1 & a_isPut & _bundleIn_0_a_ready_T_1; // @[ToAXI4.scala 199:54]
  assign deq_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_strb = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_last = counter == 3'h1 | beats1 == 3'h0; // @[Edges.scala 231:37]
  assign deq_io_deq_ready = auto_out_w_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign queue_arw_deq_clock = clock;
  assign queue_arw_deq_reset = reset;
  assign queue_arw_deq_io_enq_valid = _bundleIn_0_a_ready_T & auto_in_a_valid & _out_arw_valid_T_4; // @[ToAXI4.scala 197:45]
  assign queue_arw_deq_io_enq_bits_id = 9'h1ff == auto_in_a_bits_source ? 9'h1ff : _GEN_512; // @[ToAXI4.scala 166:{17,17}]
  assign queue_arw_deq_io_enq_bits_addr = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign queue_arw_deq_io_enq_bits_len = _out_arw_bits_len_T_3[10:3]; // @[ToAXI4.scala 168:84]
  assign queue_arw_deq_io_enq_bits_size = auto_in_a_bits_size >= 3'h3 ? 3'h3 : auto_in_a_bits_size; // @[ToAXI4.scala 169:23]
  assign queue_arw_deq_io_enq_bits_cache = {out_arw_bits_cache_hi,out_arw_bits_cache_lo}; // @[Cat.scala 31:58]
  assign queue_arw_deq_io_enq_bits_prot = {out_arw_bits_prot_hi,auto_in_a_bits_user_amba_prot_privileged}; // @[Cat.scala 31:58]
  assign queue_arw_deq_io_enq_bits_echo_tl_state_size = {{1'd0}, auto_in_a_bits_size}; // @[ToAXI4.scala 147:25 179:22]
  assign queue_arw_deq_io_enq_bits_echo_tl_state_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign queue_arw_deq_io_enq_bits_wen = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  assign queue_arw_deq_io_deq_ready = queue_arw_bits_wen ? auto_out_aw_ready : auto_out_ar_ready; // @[ToAXI4.scala 157:29]
  assign TLToAXI4_covMap_read_en = 1'h1;
  assign TLToAXI4_covMap_read_addr = TLToAXI4_covState;
  assign TLToAXI4_covMap_read_data = TLToAXI4_covMap[TLToAXI4_covMap_read_addr]; // @[Coverage map for TLToAXI4]
  assign TLToAXI4_covMap_write_data = 1'h1;
  assign TLToAXI4_covMap_write_addr = TLToAXI4_covState;
  assign TLToAXI4_covMap_write_mask = 1'h1;
  assign TLToAXI4_covMap_write_en = ~metaReset;
  assign count_331_shl = {count_331, 10'h0};
  assign count_331_pad = {9'h0,count_331_shl};
  assign count_401_shl = {count_401, 17'h0};
  assign count_401_pad = {2'h0,count_401_shl};
  assign count_227_shl = {count_227, 18'h0};
  assign count_227_pad = {1'h0,count_227_shl};
  assign count_383_shl = {count_383, 2'h0};
  assign count_383_pad = {17'h0,count_383_shl};
  assign count_195_shl = {count_195, 7'h0};
  assign count_195_pad = {12'h0,count_195_shl};
  assign count_417_shl = {count_417, 18'h0};
  assign count_417_pad = {1'h0,count_417_shl};
  assign count_121_shl = {count_121, 10'h0};
  assign count_121_pad = {9'h0,count_121_shl};
  assign count_447_shl = {count_447, 12'h0};
  assign count_447_pad = {7'h0,count_447_shl};
  assign count_482_shl = {count_482, 12'h0};
  assign count_482_pad = {7'h0,count_482_shl};
  assign count_26_shl = count_26;
  assign count_26_pad = {19'h0,count_26_shl};
  assign count_391_shl = {count_391, 17'h0};
  assign count_391_pad = {2'h0,count_391_shl};
  assign count_284_shl = {count_284, 18'h0};
  assign count_284_pad = {1'h0,count_284_shl};
  assign count_204_shl = {count_204, 4'h0};
  assign count_204_pad = {15'h0,count_204_shl};
  assign count_199_shl = {count_199, 13'h0};
  assign count_199_pad = {6'h0,count_199_shl};
  assign count_373_shl = {count_373, 4'h0};
  assign count_373_pad = {15'h0,count_373_shl};
  assign count_394_shl = {count_394, 9'h0};
  assign count_394_pad = {10'h0,count_394_shl};
  assign count_411_shl = {count_411, 13'h0};
  assign count_411_pad = {6'h0,count_411_shl};
  assign count_120_shl = {count_120, 16'h0};
  assign count_120_pad = {3'h0,count_120_shl};
  assign count_503_shl = {count_503, 17'h0};
  assign count_503_pad = {2'h0,count_503_shl};
  assign count_70_shl = {count_70, 3'h0};
  assign count_70_pad = {16'h0,count_70_shl};
  assign count_270_shl = {count_270, 8'h0};
  assign count_270_pad = {11'h0,count_270_shl};
  assign count_372_shl = {count_372, 14'h0};
  assign count_372_pad = {5'h0,count_372_shl};
  assign count_474_shl = {count_474, 12'h0};
  assign count_474_pad = {7'h0,count_474_shl};
  assign count_421_shl = {count_421, 17'h0};
  assign count_421_pad = {2'h0,count_421_shl};
  assign count_501_shl = {count_501, 6'h0};
  assign count_501_pad = {13'h0,count_501_shl};
  assign count_154_shl = {count_154, 2'h0};
  assign count_154_pad = {17'h0,count_154_shl};
  assign count_329_shl = {count_329, 9'h0};
  assign count_329_pad = {10'h0,count_329_shl};
  assign count_117_shl = {count_117, 3'h0};
  assign count_117_pad = {16'h0,count_117_shl};
  assign count_297_shl = {count_297, 12'h0};
  assign count_297_pad = {7'h0,count_297_shl};
  assign count_202_shl = {count_202, 4'h0};
  assign count_202_pad = {15'h0,count_202_shl};
  assign count_50_shl = {count_50, 5'h0};
  assign count_50_pad = {14'h0,count_50_shl};
  assign count_184_shl = {count_184, 11'h0};
  assign count_184_pad = {8'h0,count_184_shl};
  assign count_263_shl = {count_263, 7'h0};
  assign count_263_pad = {12'h0,count_263_shl};
  assign count_313_shl = {count_313, 19'h0};
  assign count_313_pad = count_313_shl;
  assign count_168_shl = {count_168, 12'h0};
  assign count_168_pad = {7'h0,count_168_shl};
  assign count_305_shl = {count_305, 2'h0};
  assign count_305_pad = {17'h0,count_305_shl};
  assign count_38_shl = {count_38, 1'h0};
  assign count_38_pad = {18'h0,count_38_shl};
  assign count_310_shl = {count_310, 1'h0};
  assign count_310_pad = {18'h0,count_310_shl};
  assign count_317_shl = {count_317, 16'h0};
  assign count_317_pad = {3'h0,count_317_shl};
  assign count_393_shl = count_393;
  assign count_393_pad = {19'h0,count_393_shl};
  assign count_182_shl = {count_182, 8'h0};
  assign count_182_pad = {11'h0,count_182_shl};
  assign count_357_shl = {count_357, 12'h0};
  assign count_357_pad = {7'h0,count_357_shl};
  assign count_423_shl = {count_423, 15'h0};
  assign count_423_pad = {4'h0,count_423_shl};
  assign count_37_shl = {count_37, 19'h0};
  assign count_37_pad = count_37_shl;
  assign count_31_shl = {count_31, 4'h0};
  assign count_31_pad = {15'h0,count_31_shl};
  assign count_61_shl = {count_61, 6'h0};
  assign count_61_pad = {13'h0,count_61_shl};
  assign count_333_shl = {count_333, 15'h0};
  assign count_333_pad = {4'h0,count_333_shl};
  assign count_296_shl = count_296;
  assign count_296_pad = {19'h0,count_296_shl};
  assign count_222_shl = {count_222, 13'h0};
  assign count_222_pad = {6'h0,count_222_shl};
  assign count_477_shl = {count_477, 17'h0};
  assign count_477_pad = {2'h0,count_477_shl};
  assign count_498_shl = {count_498, 14'h0};
  assign count_498_pad = {5'h0,count_498_shl};
  assign count_422_shl = {count_422, 10'h0};
  assign count_422_pad = {9'h0,count_422_shl};
  assign count_67_shl = {count_67, 3'h0};
  assign count_67_pad = {16'h0,count_67_shl};
  assign count_420_shl = {count_420, 1'h0};
  assign count_420_pad = {18'h0,count_420_shl};
  assign count_293_shl = {count_293, 2'h0};
  assign count_293_pad = {17'h0,count_293_shl};
  assign count_242_shl = {count_242, 15'h0};
  assign count_242_pad = {4'h0,count_242_shl};
  assign count_64_shl = {count_64, 1'h0};
  assign count_64_pad = {18'h0,count_64_shl};
  assign count_223_shl = {count_223, 7'h0};
  assign count_223_pad = {12'h0,count_223_shl};
  assign count_352_shl = {count_352, 19'h0};
  assign count_352_pad = count_352_shl;
  assign count_153_shl = {count_153, 9'h0};
  assign count_153_pad = {10'h0,count_153_shl};
  assign count_118_shl = {count_118, 14'h0};
  assign count_118_pad = {5'h0,count_118_shl};
  assign count_139_shl = {count_139, 1'h0};
  assign count_139_pad = {18'h0,count_139_shl};
  assign count_467_shl = {count_467, 8'h0};
  assign count_467_pad = {11'h0,count_467_shl};
  assign count_386_shl = {count_386, 2'h0};
  assign count_386_pad = {17'h0,count_386_shl};
  assign count_434_shl = {count_434, 6'h0};
  assign count_434_pad = {13'h0,count_434_shl};
  assign count_51_shl = {count_51, 16'h0};
  assign count_51_pad = {3'h0,count_51_shl};
  assign count_129_shl = {count_129, 13'h0};
  assign count_129_pad = {6'h0,count_129_shl};
  assign count_378_shl = {count_378, 5'h0};
  assign count_378_pad = {14'h0,count_378_shl};
  assign count_186_shl = {count_186, 10'h0};
  assign count_186_pad = {9'h0,count_186_shl};
  assign count_101_shl = {count_101, 9'h0};
  assign count_101_pad = {10'h0,count_101_shl};
  assign count_229_shl = {count_229, 19'h0};
  assign count_229_pad = count_229_shl;
  assign count_280_shl = {count_280, 10'h0};
  assign count_280_pad = {9'h0,count_280_shl};
  assign count_403_shl = {count_403, 11'h0};
  assign count_403_pad = {8'h0,count_403_shl};
  assign count_330_shl = {count_330, 8'h0};
  assign count_330_pad = {11'h0,count_330_shl};
  assign count_398_shl = {count_398, 10'h0};
  assign count_398_pad = {9'h0,count_398_shl};
  assign count_307_shl = {count_307, 4'h0};
  assign count_307_pad = {15'h0,count_307_shl};
  assign count_216_shl = {count_216, 1'h0};
  assign count_216_pad = {18'h0,count_216_shl};
  assign count_400_shl = {count_400, 6'h0};
  assign count_400_pad = {13'h0,count_400_shl};
  assign count_304_shl = {count_304, 3'h0};
  assign count_304_pad = {16'h0,count_304_shl};
  assign count_131_shl = {count_131, 13'h0};
  assign count_131_pad = {6'h0,count_131_shl};
  assign count_282_shl = {count_282, 9'h0};
  assign count_282_pad = {10'h0,count_282_shl};
  assign count_35_shl = {count_35, 11'h0};
  assign count_35_pad = {8'h0,count_35_shl};
  assign count_428_shl = {count_428, 10'h0};
  assign count_428_pad = {9'h0,count_428_shl};
  assign count_16_shl = {count_16, 14'h0};
  assign count_16_pad = {5'h0,count_16_shl};
  assign count_355_shl = {count_355, 11'h0};
  assign count_355_pad = {8'h0,count_355_shl};
  assign count_110_shl = count_110;
  assign count_110_pad = {19'h0,count_110_shl};
  assign count_367_shl = {count_367, 18'h0};
  assign count_367_pad = {1'h0,count_367_shl};
  assign count_427_shl = {count_427, 17'h0};
  assign count_427_pad = {2'h0,count_427_shl};
  assign count_46_shl = {count_46, 2'h0};
  assign count_46_pad = {17'h0,count_46_shl};
  assign count_272_shl = {count_272, 3'h0};
  assign count_272_pad = {16'h0,count_272_shl};
  assign count_5_shl = {count_5, 17'h0};
  assign count_5_pad = {2'h0,count_5_shl};
  assign count_173_shl = {count_173, 6'h0};
  assign count_173_pad = {13'h0,count_173_shl};
  assign count_211_shl = {count_211, 18'h0};
  assign count_211_pad = {1'h0,count_211_shl};
  assign count_230_shl = {count_230, 1'h0};
  assign count_230_pad = {18'h0,count_230_shl};
  assign count_454_shl = {count_454, 7'h0};
  assign count_454_pad = {12'h0,count_454_shl};
  assign count_458_shl = {count_458, 10'h0};
  assign count_458_pad = {9'h0,count_458_shl};
  assign count_23_shl = {count_23, 5'h0};
  assign count_23_pad = {14'h0,count_23_shl};
  assign count_350_shl = {count_350, 12'h0};
  assign count_350_pad = {7'h0,count_350_shl};
  assign count_368_shl = {count_368, 7'h0};
  assign count_368_pad = {12'h0,count_368_shl};
  assign count_456_shl = {count_456, 7'h0};
  assign count_456_pad = {12'h0,count_456_shl};
  assign count_464_shl = {count_464, 6'h0};
  assign count_464_pad = {13'h0,count_464_shl};
  assign count_56_shl = {count_56, 3'h0};
  assign count_56_pad = {16'h0,count_56_shl};
  assign count_158_shl = {count_158, 6'h0};
  assign count_158_pad = {13'h0,count_158_shl};
  assign count_1_shl = {count_1, 13'h0};
  assign count_1_pad = {6'h0,count_1_shl};
  assign count_62_shl = {count_62, 7'h0};
  assign count_62_pad = {12'h0,count_62_shl};
  assign count_295_shl = {count_295, 4'h0};
  assign count_295_pad = {15'h0,count_295_shl};
  assign count_285_shl = {count_285, 7'h0};
  assign count_285_pad = {12'h0,count_285_shl};
  assign count_44_shl = {count_44, 9'h0};
  assign count_44_pad = {10'h0,count_44_shl};
  assign count_25_shl = {count_25, 17'h0};
  assign count_25_pad = {2'h0,count_25_shl};
  assign count_256_shl = {count_256, 1'h0};
  assign count_256_pad = {18'h0,count_256_shl};
  assign count_366_shl = {count_366, 17'h0};
  assign count_366_pad = {2'h0,count_366_shl};
  assign count_473_shl = {count_473, 13'h0};
  assign count_473_pad = {6'h0,count_473_shl};
  assign count_465_shl = {count_465, 2'h0};
  assign count_465_pad = {17'h0,count_465_shl};
  assign count_268_shl = {count_268, 10'h0};
  assign count_268_pad = {9'h0,count_268_shl};
  assign count_142_shl = {count_142, 19'h0};
  assign count_142_pad = count_142_shl;
  assign count_75_shl = {count_75, 4'h0};
  assign count_75_pad = {15'h0,count_75_shl};
  assign count_240_shl = {count_240, 9'h0};
  assign count_240_pad = {10'h0,count_240_shl};
  assign count_481_shl = {count_481, 2'h0};
  assign count_481_pad = {17'h0,count_481_shl};
  assign count_189_shl = {count_189, 1'h0};
  assign count_189_pad = {18'h0,count_189_shl};
  assign count_382_shl = {count_382, 4'h0};
  assign count_382_pad = {15'h0,count_382_shl};
  assign count_219_shl = {count_219, 1'h0};
  assign count_219_pad = {18'h0,count_219_shl};
  assign count_365_shl = count_365;
  assign count_365_pad = {19'h0,count_365_shl};
  assign count_300_shl = {count_300, 9'h0};
  assign count_300_pad = {10'h0,count_300_shl};
  assign count_53_shl = {count_53, 13'h0};
  assign count_53_pad = {6'h0,count_53_shl};
  assign count_490_shl = {count_490, 16'h0};
  assign count_490_pad = {3'h0,count_490_shl};
  assign count_190_shl = {count_190, 19'h0};
  assign count_190_pad = count_190_shl;
  assign count_332_shl = {count_332, 9'h0};
  assign count_332_pad = {10'h0,count_332_shl};
  assign count_258_shl = {count_258, 4'h0};
  assign count_258_pad = {15'h0,count_258_shl};
  assign count_356_shl = {count_356, 18'h0};
  assign count_356_pad = {1'h0,count_356_shl};
  assign count_410_shl = {count_410, 7'h0};
  assign count_410_pad = {12'h0,count_410_shl};
  assign count_68_shl = {count_68, 5'h0};
  assign count_68_pad = {14'h0,count_68_shl};
  assign count_444_shl = {count_444, 9'h0};
  assign count_444_pad = {10'h0,count_444_shl};
  assign count_446_shl = {count_446, 14'h0};
  assign count_446_pad = {5'h0,count_446_shl};
  assign count_493_shl = {count_493, 11'h0};
  assign count_493_pad = {8'h0,count_493_shl};
  assign count_404_shl = {count_404, 5'h0};
  assign count_404_pad = {14'h0,count_404_shl};
  assign count_40_shl = {count_40, 15'h0};
  assign count_40_pad = {4'h0,count_40_shl};
  assign count_495_shl = {count_495, 14'h0};
  assign count_495_pad = {5'h0,count_495_shl};
  assign count_325_shl = {count_325, 16'h0};
  assign count_325_pad = {3'h0,count_325_shl};
  assign count_58_shl = count_58;
  assign count_58_pad = {19'h0,count_58_shl};
  assign count_201_shl = {count_201, 19'h0};
  assign count_201_pad = count_201_shl;
  assign count_107_shl = {count_107, 18'h0};
  assign count_107_pad = {1'h0,count_107_shl};
  assign count_292_shl = {count_292, 6'h0};
  assign count_292_pad = {13'h0,count_292_shl};
  assign count_462_shl = {count_462, 4'h0};
  assign count_462_pad = {15'h0,count_462_shl};
  assign count_380_shl = count_380;
  assign count_380_pad = {19'h0,count_380_shl};
  assign count_57_shl = {count_57, 16'h0};
  assign count_57_pad = {3'h0,count_57_shl};
  assign count_395_shl = {count_395, 6'h0};
  assign count_395_pad = {13'h0,count_395_shl};
  assign count_20_shl = {count_20, 18'h0};
  assign count_20_pad = {1'h0,count_20_shl};
  assign count_99_shl = {count_99, 10'h0};
  assign count_99_pad = {9'h0,count_99_shl};
  assign count_327_shl = {count_327, 19'h0};
  assign count_327_pad = count_327_shl;
  assign count_30_shl = {count_30, 1'h0};
  assign count_30_pad = {18'h0,count_30_shl};
  assign count_302_shl = {count_302, 7'h0};
  assign count_302_pad = {12'h0,count_302_shl};
  assign count_77_shl = {count_77, 14'h0};
  assign count_77_pad = {5'h0,count_77_shl};
  assign count_439_shl = {count_439, 6'h0};
  assign count_439_pad = {13'h0,count_439_shl};
  assign count_409_shl = count_409;
  assign count_409_pad = {19'h0,count_409_shl};
  assign count_443_shl = {count_443, 8'h0};
  assign count_443_pad = {11'h0,count_443_shl};
  assign count_143_shl = {count_143, 10'h0};
  assign count_143_pad = {9'h0,count_143_shl};
  assign count_165_shl = {count_165, 5'h0};
  assign count_165_pad = {14'h0,count_165_shl};
  assign count_81_shl = {count_81, 17'h0};
  assign count_81_pad = {2'h0,count_81_shl};
  assign count_346_shl = {count_346, 19'h0};
  assign count_346_pad = count_346_shl;
  assign count_314_shl = {count_314, 6'h0};
  assign count_314_pad = {13'h0,count_314_shl};
  assign count_196_shl = {count_196, 5'h0};
  assign count_196_pad = {14'h0,count_196_shl};
  assign count_262_shl = {count_262, 2'h0};
  assign count_262_pad = {17'h0,count_262_shl};
  assign count_402_shl = {count_402, 14'h0};
  assign count_402_pad = {5'h0,count_402_shl};
  assign count_87_shl = {count_87, 18'h0};
  assign count_87_pad = {1'h0,count_87_shl};
  assign count_29_shl = {count_29, 5'h0};
  assign count_29_pad = {14'h0,count_29_shl};
  assign count_126_shl = {count_126, 13'h0};
  assign count_126_pad = {6'h0,count_126_shl};
  assign count_318_shl = {count_318, 6'h0};
  assign count_318_pad = {13'h0,count_318_shl};
  assign count_66_shl = {count_66, 2'h0};
  assign count_66_pad = {17'h0,count_66_shl};
  assign count_163_shl = {count_163, 1'h0};
  assign count_163_pad = {18'h0,count_163_shl};
  assign count_175_shl = {count_175, 4'h0};
  assign count_175_pad = {15'h0,count_175_shl};
  assign count_71_shl = {count_71, 14'h0};
  assign count_71_pad = {5'h0,count_71_shl};
  assign count_80_shl = {count_80, 9'h0};
  assign count_80_pad = {10'h0,count_80_shl};
  assign count_252_shl = count_252;
  assign count_252_pad = {19'h0,count_252_shl};
  assign count_28_shl = {count_28, 6'h0};
  assign count_28_pad = {13'h0,count_28_shl};
  assign count_502_shl = {count_502, 17'h0};
  assign count_502_pad = {2'h0,count_502_shl};
  assign count_459_shl = {count_459, 19'h0};
  assign count_459_pad = count_459_shl;
  assign count_141_shl = {count_141, 15'h0};
  assign count_141_pad = {4'h0,count_141_shl};
  assign count_405_shl = {count_405, 16'h0};
  assign count_405_pad = {3'h0,count_405_shl};
  assign count_511_shl = {count_511, 3'h0};
  assign count_511_pad = {16'h0,count_511_shl};
  assign count_254_shl = {count_254, 7'h0};
  assign count_254_pad = {12'h0,count_254_shl};
  assign count_476_shl = {count_476, 15'h0};
  assign count_476_pad = {4'h0,count_476_shl};
  assign count_97_shl = {count_97, 2'h0};
  assign count_97_pad = {17'h0,count_97_shl};
  assign count_448_shl = {count_448, 3'h0};
  assign count_448_pad = {16'h0,count_448_shl};
  assign count_193_shl = {count_193, 12'h0};
  assign count_193_pad = {7'h0,count_193_shl};
  assign count_260_shl = {count_260, 16'h0};
  assign count_260_pad = {3'h0,count_260_shl};
  assign count_303_shl = {count_303, 18'h0};
  assign count_303_pad = {1'h0,count_303_shl};
  assign count_177_shl = {count_177, 6'h0};
  assign count_177_pad = {13'h0,count_177_shl};
  assign count_470_shl = {count_470, 6'h0};
  assign count_470_pad = {13'h0,count_470_shl};
  assign count_146_shl = {count_146, 8'h0};
  assign count_146_pad = {11'h0,count_146_shl};
  assign count_309_shl = count_309;
  assign count_309_pad = {19'h0,count_309_shl};
  assign count_213_shl = {count_213, 12'h0};
  assign count_213_pad = {7'h0,count_213_shl};
  assign count_343_shl = {count_343, 17'h0};
  assign count_343_pad = {2'h0,count_343_shl};
  assign count_468_shl = {count_468, 16'h0};
  assign count_468_pad = {3'h0,count_468_shl};
  assign count_429_shl = {count_429, 7'h0};
  assign count_429_pad = {12'h0,count_429_shl};
  assign count_244_shl = {count_244, 12'h0};
  assign count_244_pad = {7'h0,count_244_shl};
  assign count_69_shl = {count_69, 19'h0};
  assign count_69_pad = count_69_shl;
  assign count_460_shl = {count_460, 19'h0};
  assign count_460_pad = count_460_shl;
  assign count_370_shl = count_370;
  assign count_370_pad = {19'h0,count_370_shl};
  assign count_125_shl = {count_125, 10'h0};
  assign count_125_pad = {9'h0,count_125_shl};
  assign count_290_shl = {count_290, 12'h0};
  assign count_290_pad = {7'h0,count_290_shl};
  assign count_128_shl = count_128;
  assign count_128_pad = {19'h0,count_128_shl};
  assign count_407_shl = {count_407, 13'h0};
  assign count_407_pad = {6'h0,count_407_shl};
  assign count_198_shl = {count_198, 9'h0};
  assign count_198_pad = {10'h0,count_198_shl};
  assign count_140_shl = {count_140, 4'h0};
  assign count_140_pad = {15'h0,count_140_shl};
  assign count_512_shl = {count_512, 9'h0};
  assign count_512_pad = {10'h0,count_512_shl};
  assign count_440_shl = {count_440, 9'h0};
  assign count_440_pad = {10'h0,count_440_shl};
  assign count_362_shl = {count_362, 4'h0};
  assign count_362_pad = {15'h0,count_362_shl};
  assign count_480_shl = {count_480, 12'h0};
  assign count_480_pad = {7'h0,count_480_shl};
  assign count_109_shl = {count_109, 10'h0};
  assign count_109_pad = {9'h0,count_109_shl};
  assign count_171_shl = {count_171, 10'h0};
  assign count_171_pad = {9'h0,count_171_shl};
  assign count_414_shl = {count_414, 18'h0};
  assign count_414_pad = {1'h0,count_414_shl};
  assign count_267_shl = {count_267, 17'h0};
  assign count_267_pad = {2'h0,count_267_shl};
  assign count_484_shl = {count_484, 13'h0};
  assign count_484_pad = {6'h0,count_484_shl};
  assign count_278_shl = {count_278, 8'h0};
  assign count_278_pad = {11'h0,count_278_shl};
  assign count_39_shl = {count_39, 9'h0};
  assign count_39_pad = {10'h0,count_39_shl};
  assign count_360_shl = {count_360, 9'h0};
  assign count_360_pad = {10'h0,count_360_shl};
  assign count_14_shl = {count_14, 1'h0};
  assign count_14_pad = {18'h0,count_14_shl};
  assign count_336_shl = {count_336, 10'h0};
  assign count_336_pad = {9'h0,count_336_shl};
  assign count_108_shl = {count_108, 8'h0};
  assign count_108_pad = {11'h0,count_108_shl};
  assign count_45_shl = {count_45, 8'h0};
  assign count_45_pad = {11'h0,count_45_shl};
  assign count_275_shl = {count_275, 5'h0};
  assign count_275_pad = {14'h0,count_275_shl};
  assign count_413_shl = {count_413, 7'h0};
  assign count_413_pad = {12'h0,count_413_shl};
  assign count_52_shl = {count_52, 9'h0};
  assign count_52_pad = {10'h0,count_52_shl};
  assign count_41_shl = {count_41, 9'h0};
  assign count_41_pad = {10'h0,count_41_shl};
  assign count_328_shl = {count_328, 13'h0};
  assign count_328_pad = {6'h0,count_328_shl};
  assign count_82_shl = {count_82, 16'h0};
  assign count_82_pad = {3'h0,count_82_shl};
  assign count_4_shl = {count_4, 18'h0};
  assign count_4_pad = {1'h0,count_4_shl};
  assign count_299_shl = {count_299, 19'h0};
  assign count_299_pad = count_299_shl;
  assign count_286_shl = {count_286, 1'h0};
  assign count_286_pad = {18'h0,count_286_shl};
  assign count_510_shl = {count_510, 1'h0};
  assign count_510_pad = {18'h0,count_510_shl};
  assign count_96_shl = {count_96, 11'h0};
  assign count_96_pad = {8'h0,count_96_shl};
  assign count_203_shl = {count_203, 7'h0};
  assign count_203_pad = {12'h0,count_203_shl};
  assign count_452_shl = {count_452, 15'h0};
  assign count_452_pad = {4'h0,count_452_shl};
  assign count_150_shl = {count_150, 13'h0};
  assign count_150_pad = {6'h0,count_150_shl};
  assign count_385_shl = {count_385, 2'h0};
  assign count_385_pad = {17'h0,count_385_shl};
  assign count_156_shl = {count_156, 7'h0};
  assign count_156_pad = {12'h0,count_156_shl};
  assign count_169_shl = {count_169, 15'h0};
  assign count_169_pad = {4'h0,count_169_shl};
  assign count_132_shl = {count_132, 10'h0};
  assign count_132_pad = {9'h0,count_132_shl};
  assign count_225_shl = {count_225, 12'h0};
  assign count_225_pad = {7'h0,count_225_shl};
  assign count_341_shl = {count_341, 19'h0};
  assign count_341_pad = count_341_shl;
  assign count_377_shl = {count_377, 2'h0};
  assign count_377_pad = {17'h0,count_377_shl};
  assign count_114_shl = {count_114, 6'h0};
  assign count_114_pad = {13'h0,count_114_shl};
  assign count_294_shl = {count_294, 7'h0};
  assign count_294_pad = {12'h0,count_294_shl};
  assign count_79_shl = {count_79, 12'h0};
  assign count_79_pad = {7'h0,count_79_shl};
  assign count_60_shl = {count_60, 15'h0};
  assign count_60_pad = {4'h0,count_60_shl};
  assign count_86_shl = {count_86, 1'h0};
  assign count_86_pad = {18'h0,count_86_shl};
  assign count_399_shl = {count_399, 14'h0};
  assign count_399_pad = {5'h0,count_399_shl};
  assign count_279_shl = {count_279, 15'h0};
  assign count_279_pad = {4'h0,count_279_shl};
  assign count_239_shl = {count_239, 15'h0};
  assign count_239_pad = {4'h0,count_239_shl};
  assign count_13_shl = {count_13, 12'h0};
  assign count_13_pad = {7'h0,count_13_shl};
  assign count_337_shl = {count_337, 16'h0};
  assign count_337_pad = {3'h0,count_337_shl};
  assign count_19_shl = {count_19, 5'h0};
  assign count_19_pad = {14'h0,count_19_shl};
  assign count_334_shl = {count_334, 9'h0};
  assign count_334_pad = {10'h0,count_334_shl};
  assign count_17_shl = {count_17, 16'h0};
  assign count_17_pad = {3'h0,count_17_shl};
  assign count_72_shl = {count_72, 5'h0};
  assign count_72_pad = {14'h0,count_72_shl};
  assign count_94_shl = {count_94, 14'h0};
  assign count_94_pad = {5'h0,count_94_shl};
  assign count_419_shl = {count_419, 5'h0};
  assign count_419_pad = {14'h0,count_419_shl};
  assign count_176_shl = count_176;
  assign count_176_pad = {19'h0,count_176_shl};
  assign count_210_shl = {count_210, 11'h0};
  assign count_210_pad = {8'h0,count_210_shl};
  assign count_78_shl = {count_78, 14'h0};
  assign count_78_pad = {5'h0,count_78_shl};
  assign count_104_shl = {count_104, 17'h0};
  assign count_104_pad = {2'h0,count_104_shl};
  assign count_507_shl = {count_507, 19'h0};
  assign count_507_pad = count_507_shl;
  assign count_287_shl = {count_287, 17'h0};
  assign count_287_pad = {2'h0,count_287_shl};
  assign count_208_shl = count_208;
  assign count_208_pad = {19'h0,count_208_shl};
  assign count_345_shl = {count_345, 9'h0};
  assign count_345_pad = {10'h0,count_345_shl};
  assign count_311_shl = {count_311, 14'h0};
  assign count_311_pad = {5'h0,count_311_shl};
  assign count_178_shl = {count_178, 3'h0};
  assign count_178_pad = {16'h0,count_178_shl};
  assign count_89_shl = {count_89, 6'h0};
  assign count_89_pad = {13'h0,count_89_shl};
  assign count_266_shl = {count_266, 17'h0};
  assign count_266_pad = {2'h0,count_266_shl};
  assign count_238_shl = {count_238, 2'h0};
  assign count_238_pad = {17'h0,count_238_shl};
  assign count_206_shl = {count_206, 5'h0};
  assign count_206_pad = {14'h0,count_206_shl};
  assign count_103_shl = {count_103, 18'h0};
  assign count_103_pad = {1'h0,count_103_shl};
  assign count_85_shl = {count_85, 15'h0};
  assign count_85_pad = {4'h0,count_85_shl};
  assign count_138_shl = {count_138, 15'h0};
  assign count_138_pad = {4'h0,count_138_shl};
  assign count_392_shl = {count_392, 18'h0};
  assign count_392_pad = {1'h0,count_392_shl};
  assign count_271_shl = {count_271, 16'h0};
  assign count_271_pad = {3'h0,count_271_shl};
  assign count_445_shl = {count_445, 15'h0};
  assign count_445_pad = {4'h0,count_445_shl};
  assign count_431_shl = {count_431, 10'h0};
  assign count_431_pad = {9'h0,count_431_shl};
  assign count_220_shl = {count_220, 14'h0};
  assign count_220_pad = {5'h0,count_220_shl};
  assign count_160_shl = {count_160, 9'h0};
  assign count_160_pad = {10'h0,count_160_shl};
  assign count_183_shl = {count_183, 11'h0};
  assign count_183_pad = {8'h0,count_183_shl};
  assign count_436_shl = {count_436, 13'h0};
  assign count_436_pad = {6'h0,count_436_shl};
  assign count_226_shl = {count_226, 19'h0};
  assign count_226_pad = count_226_shl;
  assign count_136_shl = {count_136, 16'h0};
  assign count_136_pad = {3'h0,count_136_shl};
  assign count_42_shl = {count_42, 18'h0};
  assign count_42_pad = {1'h0,count_42_shl};
  assign count_351_shl = count_351;
  assign count_351_pad = {19'h0,count_351_shl};
  assign count_261_shl = {count_261, 17'h0};
  assign count_261_pad = {2'h0,count_261_shl};
  assign count_221_shl = {count_221, 4'h0};
  assign count_221_pad = {15'h0,count_221_shl};
  assign count_152_shl = count_152;
  assign count_152_pad = {19'h0,count_152_shl};
  assign count_505_shl = {count_505, 7'h0};
  assign count_505_pad = {12'h0,count_505_shl};
  assign count_36_shl = {count_36, 9'h0};
  assign count_36_pad = {10'h0,count_36_shl};
  assign count_232_shl = {count_232, 13'h0};
  assign count_232_pad = {6'h0,count_232_shl};
  assign count_479_shl = {count_479, 5'h0};
  assign count_479_pad = {14'h0,count_479_shl};
  assign count_34_shl = {count_34, 19'h0};
  assign count_34_pad = count_34_shl;
  assign count_291_shl = {count_291, 4'h0};
  assign count_291_pad = {15'h0,count_291_shl};
  assign count_246_shl = {count_246, 11'h0};
  assign count_246_pad = {8'h0,count_246_shl};
  assign count_9_shl = {count_9, 15'h0};
  assign count_9_pad = {4'h0,count_9_shl};
  assign count_98_shl = {count_98, 3'h0};
  assign count_98_pad = {16'h0,count_98_shl};
  assign count_364_shl = {count_364, 1'h0};
  assign count_364_pad = {18'h0,count_364_shl};
  assign count_451_shl = {count_451, 14'h0};
  assign count_451_pad = {5'h0,count_451_shl};
  assign count_426_shl = {count_426, 16'h0};
  assign count_426_pad = {3'h0,count_426_shl};
  assign count_492_shl = {count_492, 1'h0};
  assign count_492_pad = {18'h0,count_492_shl};
  assign count_281_shl = {count_281, 4'h0};
  assign count_281_pad = {15'h0,count_281_shl};
  assign count_494_shl = count_494;
  assign count_494_pad = {19'h0,count_494_shl};
  assign count_340_shl = {count_340, 13'h0};
  assign count_340_pad = {6'h0,count_340_shl};
  assign count_179_shl = {count_179, 9'h0};
  assign count_179_pad = {10'h0,count_179_shl};
  assign count_250_shl = {count_250, 16'h0};
  assign count_250_pad = {3'h0,count_250_shl};
  assign count_249_shl = {count_249, 10'h0};
  assign count_249_pad = {9'h0,count_249_shl};
  assign count_59_shl = {count_59, 8'h0};
  assign count_59_pad = {11'h0,count_59_shl};
  assign count_320_shl = {count_320, 6'h0};
  assign count_320_pad = {13'h0,count_320_shl};
  assign count_321_shl = {count_321, 16'h0};
  assign count_321_pad = {3'h0,count_321_shl};
  assign count_449_shl = {count_449, 14'h0};
  assign count_449_pad = {5'h0,count_449_shl};
  assign count_2_shl = {count_2, 8'h0};
  assign count_2_pad = {11'h0,count_2_shl};
  assign count_496_shl = {count_496, 11'h0};
  assign count_496_pad = {8'h0,count_496_shl};
  assign count_188_shl = {count_188, 2'h0};
  assign count_188_pad = {17'h0,count_188_shl};
  assign count_466_shl = {count_466, 13'h0};
  assign count_466_pad = {6'h0,count_466_shl};
  assign count_212_shl = {count_212, 18'h0};
  assign count_212_pad = {1'h0,count_212_shl};
  assign count_11_shl = {count_11, 18'h0};
  assign count_11_pad = {1'h0,count_11_shl};
  assign count_55_shl = {count_55, 16'h0};
  assign count_55_pad = {3'h0,count_55_shl};
  assign count_119_shl = {count_119, 2'h0};
  assign count_119_pad = {17'h0,count_119_shl};
  assign count_149_shl = {count_149, 10'h0};
  assign count_149_pad = {9'h0,count_149_shl};
  assign count_450_shl = {count_450, 9'h0};
  assign count_450_pad = {10'h0,count_450_shl};
  assign count_32_shl = {count_32, 11'h0};
  assign count_32_pad = {8'h0,count_32_shl};
  assign count_319_shl = {count_319, 19'h0};
  assign count_319_pad = count_319_shl;
  assign count_384_shl = {count_384, 1'h0};
  assign count_384_pad = {18'h0,count_384_shl};
  assign count_162_shl = {count_162, 9'h0};
  assign count_162_pad = {10'h0,count_162_shl};
  assign count_231_shl = {count_231, 14'h0};
  assign count_231_pad = {5'h0,count_231_shl};
  assign count_63_shl = {count_63, 8'h0};
  assign count_63_pad = {11'h0,count_63_shl};
  assign count_489_shl = {count_489, 5'h0};
  assign count_489_pad = {14'h0,count_489_shl};
  assign count_509_shl = {count_509, 4'h0};
  assign count_509_pad = {15'h0,count_509_shl};
  assign count_133_shl = {count_133, 1'h0};
  assign count_133_pad = {18'h0,count_133_shl};
  assign count_415_shl = {count_415, 10'h0};
  assign count_415_pad = {9'h0,count_415_shl};
  assign count_323_shl = {count_323, 7'h0};
  assign count_323_pad = {12'h0,count_323_shl};
  assign count_289_shl = {count_289, 2'h0};
  assign count_289_pad = {17'h0,count_289_shl};
  assign count_342_shl = {count_342, 1'h0};
  assign count_342_pad = {18'h0,count_342_shl};
  assign count_408_shl = {count_408, 5'h0};
  assign count_408_pad = {14'h0,count_408_shl};
  assign count_22_shl = {count_22, 8'h0};
  assign count_22_pad = {11'h0,count_22_shl};
  assign count_308_shl = {count_308, 9'h0};
  assign count_308_pad = {10'h0,count_308_shl};
  assign count_424_shl = {count_424, 15'h0};
  assign count_424_pad = {4'h0,count_424_shl};
  assign count_353_shl = {count_353, 2'h0};
  assign count_353_pad = {17'h0,count_353_shl};
  assign count_217_shl = {count_217, 3'h0};
  assign count_217_pad = {16'h0,count_217_shl};
  assign count_497_shl = {count_497, 2'h0};
  assign count_497_pad = {17'h0,count_497_shl};
  assign count_430_shl = {count_430, 12'h0};
  assign count_430_pad = {7'h0,count_430_shl};
  assign count_369_shl = {count_369, 4'h0};
  assign count_369_pad = {15'h0,count_369_shl};
  assign count_463_shl = {count_463, 12'h0};
  assign count_463_pad = {7'h0,count_463_shl};
  assign count_389_shl = count_389;
  assign count_389_pad = {19'h0,count_389_shl};
  assign count_499_shl = {count_499, 3'h0};
  assign count_499_pad = {16'h0,count_499_shl};
  assign count_315_shl = {count_315, 13'h0};
  assign count_315_pad = {6'h0,count_315_shl};
  assign count_113_shl = {count_113, 5'h0};
  assign count_113_pad = {14'h0,count_113_shl};
  assign count_506_shl = {count_506, 12'h0};
  assign count_506_pad = {7'h0,count_506_shl};
  assign count_257_shl = {count_257, 19'h0};
  assign count_257_pad = count_257_shl;
  assign count_12_shl = {count_12, 10'h0};
  assign count_12_pad = {9'h0,count_12_shl};
  assign count_397_shl = {count_397, 18'h0};
  assign count_397_pad = {1'h0,count_397_shl};
  assign count_326_shl = {count_326, 10'h0};
  assign count_326_pad = {9'h0,count_326_shl};
  assign count_469_shl = {count_469, 13'h0};
  assign count_469_pad = {6'h0,count_469_shl};
  assign count_316_shl = {count_316, 17'h0};
  assign count_316_pad = {2'h0,count_316_shl};
  assign count_248_shl = {count_248, 11'h0};
  assign count_248_pad = {8'h0,count_248_shl};
  assign r_first_shl = {r_first, 12'h0};
  assign r_first_pad = {7'h0,r_first_shl};
  assign count_390_shl = {count_390, 18'h0};
  assign count_390_pad = {1'h0,count_390_shl};
  assign count_277_shl = {count_277, 19'h0};
  assign count_277_pad = count_277_shl;
  assign count_269_shl = {count_269, 7'h0};
  assign count_269_pad = {12'h0,count_269_shl};
  assign count_218_shl = {count_218, 10'h0};
  assign count_218_pad = {9'h0,count_218_shl};
  assign count_115_shl = {count_115, 13'h0};
  assign count_115_pad = {6'h0,count_115_shl};
  assign count_166_shl = {count_166, 14'h0};
  assign count_166_pad = {5'h0,count_166_shl};
  assign count_487_shl = {count_487, 18'h0};
  assign count_487_pad = {1'h0,count_487_shl};
  assign count_192_shl = {count_192, 2'h0};
  assign count_192_pad = {17'h0,count_192_shl};
  assign count_508_shl = {count_508, 19'h0};
  assign count_508_pad = count_508_shl;
  assign count_358_shl = {count_358, 8'h0};
  assign count_358_pad = {11'h0,count_358_shl};
  assign count_416_shl = {count_416, 15'h0};
  assign count_416_pad = {4'h0,count_416_shl};
  assign count_151_shl = {count_151, 9'h0};
  assign count_151_pad = {10'h0,count_151_shl};
  assign count_354_shl = {count_354, 12'h0};
  assign count_354_pad = {7'h0,count_354_shl};
  assign count_21_shl = {count_21, 19'h0};
  assign count_21_pad = count_21_shl;
  assign r_holds_d_shl = {r_holds_d, 18'h0};
  assign r_holds_d_pad = {1'h0,r_holds_d_shl};
  assign count_339_shl = {count_339, 18'h0};
  assign count_339_pad = {1'h0,count_339_shl};
  assign count_111_shl = {count_111, 15'h0};
  assign count_111_pad = {4'h0,count_111_shl};
  assign count_18_shl = {count_18, 17'h0};
  assign count_18_pad = {2'h0,count_18_shl};
  assign count_425_shl = {count_425, 17'h0};
  assign count_425_pad = {2'h0,count_425_shl};
  assign count_455_shl = {count_455, 19'h0};
  assign count_455_pad = count_455_shl;
  assign count_437_shl = {count_437, 4'h0};
  assign count_437_pad = {15'h0,count_437_shl};
  assign count_245_shl = {count_245, 16'h0};
  assign count_245_pad = {3'h0,count_245_shl};
  assign count_116_shl = {count_116, 10'h0};
  assign count_116_pad = {9'h0,count_116_shl};
  assign count_194_shl = {count_194, 3'h0};
  assign count_194_pad = {16'h0,count_194_shl};
  assign count_127_shl = {count_127, 5'h0};
  assign count_127_pad = {14'h0,count_127_shl};
  assign count_137_shl = {count_137, 6'h0};
  assign count_137_pad = {13'h0,count_137_shl};
  assign count_483_shl = {count_483, 2'h0};
  assign count_483_pad = {17'h0,count_483_shl};
  assign count_159_shl = {count_159, 3'h0};
  assign count_159_pad = {16'h0,count_159_shl};
  assign count_301_shl = {count_301, 15'h0};
  assign count_301_pad = {4'h0,count_301_shl};
  assign count_215_shl = {count_215, 18'h0};
  assign count_215_pad = {1'h0,count_215_shl};
  assign count_288_shl = {count_288, 9'h0};
  assign count_288_pad = {10'h0,count_288_shl};
  assign count_54_shl = {count_54, 5'h0};
  assign count_54_pad = {14'h0,count_54_shl};
  assign count_27_shl = {count_27, 18'h0};
  assign count_27_pad = {1'h0,count_27_shl};
  assign count_161_shl = {count_161, 16'h0};
  assign count_161_pad = {3'h0,count_161_shl};
  assign count_106_shl = {count_106, 1'h0};
  assign count_106_pad = {18'h0,count_106_shl};
  assign count_485_shl = {count_485, 7'h0};
  assign count_485_pad = {12'h0,count_485_shl};
  assign count_259_shl = {count_259, 3'h0};
  assign count_259_pad = {16'h0,count_259_shl};
  assign count_264_shl = {count_264, 11'h0};
  assign count_264_pad = {8'h0,count_264_shl};
  assign count_91_shl = {count_91, 9'h0};
  assign count_91_pad = {10'h0,count_91_shl};
  assign count_84_shl = {count_84, 1'h0};
  assign count_84_pad = {18'h0,count_84_shl};
  assign count_312_shl = {count_312, 3'h0};
  assign count_312_pad = {16'h0,count_312_shl};
  assign count_207_shl = {count_207, 3'h0};
  assign count_207_pad = {16'h0,count_207_shl};
  assign count_172_shl = {count_172, 7'h0};
  assign count_172_pad = {12'h0,count_172_shl};
  assign count_253_shl = {count_253, 11'h0};
  assign count_253_pad = {8'h0,count_253_shl};
  assign count_148_shl = {count_148, 12'h0};
  assign count_148_pad = {7'h0,count_148_shl};
  assign count_228_shl = {count_228, 1'h0};
  assign count_228_pad = {18'h0,count_228_shl};
  assign count_10_shl = {count_10, 3'h0};
  assign count_10_pad = {16'h0,count_10_shl};
  assign count_322_shl = {count_322, 9'h0};
  assign count_322_pad = {10'h0,count_322_shl};
  assign count_363_shl = {count_363, 9'h0};
  assign count_363_pad = {10'h0,count_363_shl};
  assign count_48_shl = {count_48, 11'h0};
  assign count_48_pad = {8'h0,count_48_shl};
  assign count_236_shl = {count_236, 16'h0};
  assign count_236_pad = {3'h0,count_236_shl};
  assign count_205_shl = {count_205, 16'h0};
  assign count_205_pad = {3'h0,count_205_shl};
  assign count_191_shl = {count_191, 15'h0};
  assign count_191_pad = {4'h0,count_191_shl};
  assign count_338_shl = {count_338, 4'h0};
  assign count_338_pad = {15'h0,count_338_shl};
  assign count_276_shl = {count_276, 16'h0};
  assign count_276_pad = {3'h0,count_276_shl};
  assign count_475_shl = {count_475, 2'h0};
  assign count_475_pad = {17'h0,count_475_shl};
  assign count_24_shl = {count_24, 15'h0};
  assign count_24_pad = {4'h0,count_24_shl};
  assign count_387_shl = {count_387, 16'h0};
  assign count_387_pad = {3'h0,count_387_shl};
  assign count_438_shl = {count_438, 8'h0};
  assign count_438_pad = {11'h0,count_438_shl};
  assign count_472_shl = {count_472, 3'h0};
  assign count_472_pad = {16'h0,count_472_shl};
  assign count_167_shl = count_167;
  assign count_167_pad = {19'h0,count_167_shl};
  assign count_233_shl = {count_233, 2'h0};
  assign count_233_pad = {17'h0,count_233_shl};
  assign count_185_shl = {count_185, 6'h0};
  assign count_185_pad = {13'h0,count_185_shl};
  assign count_135_shl = {count_135, 12'h0};
  assign count_135_pad = {7'h0,count_135_shl};
  assign count_197_shl = {count_197, 18'h0};
  assign count_197_pad = {1'h0,count_197_shl};
  assign count_273_shl = {count_273, 19'h0};
  assign count_273_pad = count_273_shl;
  assign count_441_shl = {count_441, 14'h0};
  assign count_441_pad = {5'h0,count_441_shl};
  assign count_88_shl = {count_88, 1'h0};
  assign count_88_pad = {18'h0,count_88_shl};
  assign count_471_shl = {count_471, 13'h0};
  assign count_471_pad = {6'h0,count_471_shl};
  assign count_147_shl = {count_147, 9'h0};
  assign count_147_pad = {10'h0,count_147_shl};
  assign count_412_shl = {count_412, 17'h0};
  assign count_412_pad = {2'h0,count_412_shl};
  assign count_488_shl = {count_488, 18'h0};
  assign count_488_pad = {1'h0,count_488_shl};
  assign count_486_shl = {count_486, 8'h0};
  assign count_486_pad = {11'h0,count_486_shl};
  assign count_298_shl = count_298;
  assign count_298_pad = {19'h0,count_298_shl};
  assign count_442_shl = {count_442, 8'h0};
  assign count_442_pad = {11'h0,count_442_shl};
  assign count_73_shl = {count_73, 9'h0};
  assign count_73_pad = {10'h0,count_73_shl};
  assign count_237_shl = {count_237, 13'h0};
  assign count_237_pad = {6'h0,count_237_shl};
  assign count_435_shl = {count_435, 12'h0};
  assign count_435_pad = {7'h0,count_435_shl};
  assign count_6_shl = {count_6, 6'h0};
  assign count_6_pad = {13'h0,count_6_shl};
  assign count_361_shl = count_361;
  assign count_361_pad = {19'h0,count_361_shl};
  assign count_15_shl = {count_15, 1'h0};
  assign count_15_pad = {18'h0,count_15_shl};
  assign count_388_shl = {count_388, 12'h0};
  assign count_388_pad = {7'h0,count_388_shl};
  assign count_164_shl = count_164;
  assign count_164_pad = {19'h0,count_164_shl};
  assign count_255_shl = {count_255, 3'h0};
  assign count_255_pad = {16'h0,count_255_shl};
  assign count_306_shl = {count_306, 18'h0};
  assign count_306_pad = {1'h0,count_306_shl};
  assign count_381_shl = {count_381, 19'h0};
  assign count_381_pad = count_381_shl;
  assign count_130_shl = {count_130, 6'h0};
  assign count_130_pad = {13'h0,count_130_shl};
  assign count_145_shl = {count_145, 18'h0};
  assign count_145_pad = {1'h0,count_145_shl};
  assign count_8_shl = {count_8, 5'h0};
  assign count_8_pad = {14'h0,count_8_shl};
  assign count_224_shl = {count_224, 6'h0};
  assign count_224_pad = {13'h0,count_224_shl};
  assign count_349_shl = {count_349, 12'h0};
  assign count_349_pad = {7'h0,count_349_shl};
  assign count_375_shl = {count_375, 18'h0};
  assign count_375_pad = {1'h0,count_375_shl};
  assign count_457_shl = {count_457, 18'h0};
  assign count_457_pad = {1'h0,count_457_shl};
  assign b_delay_shl = {b_delay, 6'h0};
  assign b_delay_pad = {11'h0,b_delay_shl};
  assign count_181_shl = {count_181, 15'h0};
  assign count_181_pad = {4'h0,count_181_shl};
  assign count_170_shl = {count_170, 13'h0};
  assign count_170_pad = {6'h0,count_170_shl};
  assign count_3_shl = {count_3, 7'h0};
  assign count_3_pad = {12'h0,count_3_shl};
  assign count_461_shl = count_461;
  assign count_461_pad = {19'h0,count_461_shl};
  assign count_102_shl = {count_102, 11'h0};
  assign count_102_pad = {8'h0,count_102_shl};
  assign count_134_shl = {count_134, 2'h0};
  assign count_134_pad = {17'h0,count_134_shl};
  assign count_234_shl = {count_234, 17'h0};
  assign count_234_pad = {2'h0,count_234_shl};
  assign count_335_shl = {count_335, 19'h0};
  assign count_335_pad = count_335_shl;
  assign count_95_shl = {count_95, 12'h0};
  assign count_95_pad = {7'h0,count_95_shl};
  assign count_374_shl = {count_374, 6'h0};
  assign count_374_pad = {13'h0,count_374_shl};
  assign count_49_shl = {count_49, 2'h0};
  assign count_49_pad = {17'h0,count_49_shl};
  assign count_100_shl = {count_100, 8'h0};
  assign count_100_pad = {11'h0,count_100_shl};
  assign count_283_shl = {count_283, 6'h0};
  assign count_283_pad = {13'h0,count_283_shl};
  assign count_90_shl = {count_90, 17'h0};
  assign count_90_pad = {2'h0,count_90_shl};
  assign count_155_shl = {count_155, 9'h0};
  assign count_155_pad = {10'h0,count_155_shl};
  assign count_274_shl = {count_274, 1'h0};
  assign count_274_pad = {18'h0,count_274_shl};
  assign count_83_shl = {count_83, 13'h0};
  assign count_83_pad = {6'h0,count_83_shl};
  assign count_112_shl = {count_112, 11'h0};
  assign count_112_pad = {8'h0,count_112_shl};
  assign count_433_shl = {count_433, 12'h0};
  assign count_433_pad = {7'h0,count_433_shl};
  assign count_93_shl = {count_93, 1'h0};
  assign count_93_pad = {18'h0,count_93_shl};
  assign count_65_shl = {count_65, 3'h0};
  assign count_65_pad = {16'h0,count_65_shl};
  assign count_235_shl = count_235;
  assign count_235_pad = {19'h0,count_235_shl};
  assign count_371_shl = {count_371, 3'h0};
  assign count_371_pad = {16'h0,count_371_shl};
  assign count_122_shl = {count_122, 5'h0};
  assign count_122_pad = {14'h0,count_122_shl};
  assign count_247_shl = {count_247, 13'h0};
  assign count_247_pad = {6'h0,count_247_shl};
  assign count_157_shl = {count_157, 11'h0};
  assign count_157_pad = {8'h0,count_157_shl};
  assign count_180_shl = {count_180, 6'h0};
  assign count_180_pad = {13'h0,count_180_shl};
  assign count_347_shl = {count_347, 13'h0};
  assign count_347_pad = {6'h0,count_347_shl};
  assign count_251_shl = {count_251, 16'h0};
  assign count_251_pad = {3'h0,count_251_shl};
  assign count_200_shl = {count_200, 15'h0};
  assign count_200_pad = {4'h0,count_200_shl};
  assign count_187_shl = {count_187, 8'h0};
  assign count_187_pad = {11'h0,count_187_shl};
  assign count_432_shl = {count_432, 5'h0};
  assign count_432_pad = {14'h0,count_432_shl};
  assign count_123_shl = {count_123, 2'h0};
  assign count_123_pad = {17'h0,count_123_shl};
  assign count_418_shl = {count_418, 3'h0};
  assign count_418_pad = {16'h0,count_418_shl};
  assign count_406_shl = {count_406, 4'h0};
  assign count_406_pad = {15'h0,count_406_shl};
  assign count_241_shl = {count_241, 18'h0};
  assign count_241_pad = {1'h0,count_241_shl};
  assign count_33_shl = count_33;
  assign count_33_pad = {19'h0,count_33_shl};
  assign count_324_shl = {count_324, 12'h0};
  assign count_324_pad = {7'h0,count_324_shl};
  assign count_105_shl = {count_105, 5'h0};
  assign count_105_pad = {14'h0,count_105_shl};
  assign count_92_shl = {count_92, 1'h0};
  assign count_92_pad = {18'h0,count_92_shl};
  assign count_7_shl = {count_7, 5'h0};
  assign count_7_pad = {14'h0,count_7_shl};
  assign count_214_shl = count_214;
  assign count_214_pad = {19'h0,count_214_shl};
  assign count_379_shl = {count_379, 11'h0};
  assign count_379_pad = {8'h0,count_379_shl};
  assign count_359_shl = {count_359, 7'h0};
  assign count_359_pad = {12'h0,count_359_shl};
  assign doneAW_shl = {doneAW, 16'h0};
  assign doneAW_pad = {3'h0,doneAW_shl};
  assign count_144_shl = {count_144, 6'h0};
  assign count_144_pad = {13'h0,count_144_shl};
  assign count_396_shl = {count_396, 18'h0};
  assign count_396_pad = {1'h0,count_396_shl};
  assign count_376_shl = {count_376, 4'h0};
  assign count_376_pad = {15'h0,count_376_shl};
  assign count_504_shl = {count_504, 18'h0};
  assign count_504_pad = {1'h0,count_504_shl};
  assign count_124_shl = {count_124, 6'h0};
  assign count_124_pad = {13'h0,count_124_shl};
  assign count_500_shl = {count_500, 13'h0};
  assign count_500_pad = {6'h0,count_500_shl};
  assign count_209_shl = {count_209, 18'h0};
  assign count_209_pad = {1'h0,count_209_shl};
  assign count_348_shl = {count_348, 19'h0};
  assign count_348_pad = count_348_shl;
  assign count_344_shl = {count_344, 16'h0};
  assign count_344_pad = {3'h0,count_344_shl};
  assign count_76_shl = {count_76, 16'h0};
  assign count_76_pad = {3'h0,count_76_shl};
  assign count_265_shl = {count_265, 5'h0};
  assign count_265_pad = {14'h0,count_265_shl};
  assign count_453_shl = {count_453, 7'h0};
  assign count_453_pad = {12'h0,count_453_shl};
  assign count_47_shl = {count_47, 9'h0};
  assign count_47_pad = {10'h0,count_47_shl};
  assign count_43_shl = {count_43, 2'h0};
  assign count_43_pad = {17'h0,count_43_shl};
  assign count_74_shl = {count_74, 5'h0};
  assign count_74_pad = {14'h0,count_74_shl};
  assign count_491_shl = {count_491, 6'h0};
  assign count_491_pad = {13'h0,count_491_shl};
  assign count_478_shl = {count_478, 9'h0};
  assign count_478_pad = {10'h0,count_478_shl};
  assign count_243_shl = {count_243, 6'h0};
  assign count_243_pad = {13'h0,count_243_shl};
  assign count_174_shl = count_174;
  assign count_174_pad = {19'h0,count_174_shl};
  assign TLToAXI4_xor255 = count_331_pad ^ count_401_pad;
  assign TLToAXI4_xor256 = count_227_pad ^ count_383_pad;
  assign TLToAXI4_xor127 = TLToAXI4_xor255 ^ TLToAXI4_xor256;
  assign TLToAXI4_xor257 = count_195_pad ^ count_417_pad;
  assign TLToAXI4_xor258 = count_121_pad ^ count_447_pad;
  assign TLToAXI4_xor128 = TLToAXI4_xor257 ^ TLToAXI4_xor258;
  assign TLToAXI4_xor63 = TLToAXI4_xor127 ^ TLToAXI4_xor128;
  assign TLToAXI4_xor259 = count_482_pad ^ count_26_pad;
  assign TLToAXI4_xor260 = count_391_pad ^ count_284_pad;
  assign TLToAXI4_xor129 = TLToAXI4_xor259 ^ TLToAXI4_xor260;
  assign TLToAXI4_xor261 = count_204_pad ^ count_199_pad;
  assign TLToAXI4_xor262 = count_373_pad ^ count_394_pad;
  assign TLToAXI4_xor130 = TLToAXI4_xor261 ^ TLToAXI4_xor262;
  assign TLToAXI4_xor64 = TLToAXI4_xor129 ^ TLToAXI4_xor130;
  assign TLToAXI4_xor31 = TLToAXI4_xor63 ^ TLToAXI4_xor64;
  assign TLToAXI4_xor263 = count_411_pad ^ count_120_pad;
  assign TLToAXI4_xor264 = count_503_pad ^ count_70_pad;
  assign TLToAXI4_xor131 = TLToAXI4_xor263 ^ TLToAXI4_xor264;
  assign TLToAXI4_xor265 = count_270_pad ^ count_372_pad;
  assign TLToAXI4_xor266 = count_474_pad ^ count_421_pad;
  assign TLToAXI4_xor132 = TLToAXI4_xor265 ^ TLToAXI4_xor266;
  assign TLToAXI4_xor65 = TLToAXI4_xor131 ^ TLToAXI4_xor132;
  assign TLToAXI4_xor267 = count_501_pad ^ count_154_pad;
  assign TLToAXI4_xor268 = count_329_pad ^ count_117_pad;
  assign TLToAXI4_xor133 = TLToAXI4_xor267 ^ TLToAXI4_xor268;
  assign TLToAXI4_xor269 = count_297_pad ^ count_202_pad;
  assign TLToAXI4_xor270 = count_50_pad ^ count_184_pad;
  assign TLToAXI4_xor134 = TLToAXI4_xor269 ^ TLToAXI4_xor270;
  assign TLToAXI4_xor66 = TLToAXI4_xor133 ^ TLToAXI4_xor134;
  assign TLToAXI4_xor32 = TLToAXI4_xor65 ^ TLToAXI4_xor66;
  assign TLToAXI4_xor15 = TLToAXI4_xor31 ^ TLToAXI4_xor32;
  assign TLToAXI4_xor271 = count_263_pad ^ count_313_pad;
  assign TLToAXI4_xor272 = count_168_pad ^ count_305_pad;
  assign TLToAXI4_xor135 = TLToAXI4_xor271 ^ TLToAXI4_xor272;
  assign TLToAXI4_xor273 = count_38_pad ^ count_310_pad;
  assign TLToAXI4_xor274 = count_317_pad ^ count_393_pad;
  assign TLToAXI4_xor136 = TLToAXI4_xor273 ^ TLToAXI4_xor274;
  assign TLToAXI4_xor67 = TLToAXI4_xor135 ^ TLToAXI4_xor136;
  assign TLToAXI4_xor275 = count_182_pad ^ count_357_pad;
  assign TLToAXI4_xor276 = count_423_pad ^ count_37_pad;
  assign TLToAXI4_xor137 = TLToAXI4_xor275 ^ TLToAXI4_xor276;
  assign TLToAXI4_xor277 = count_31_pad ^ count_61_pad;
  assign TLToAXI4_xor278 = count_333_pad ^ count_296_pad;
  assign TLToAXI4_xor138 = TLToAXI4_xor277 ^ TLToAXI4_xor278;
  assign TLToAXI4_xor68 = TLToAXI4_xor137 ^ TLToAXI4_xor138;
  assign TLToAXI4_xor33 = TLToAXI4_xor67 ^ TLToAXI4_xor68;
  assign TLToAXI4_xor279 = count_222_pad ^ count_477_pad;
  assign TLToAXI4_xor280 = count_498_pad ^ count_422_pad;
  assign TLToAXI4_xor139 = TLToAXI4_xor279 ^ TLToAXI4_xor280;
  assign TLToAXI4_xor281 = count_67_pad ^ count_420_pad;
  assign TLToAXI4_xor282 = count_293_pad ^ count_242_pad;
  assign TLToAXI4_xor140 = TLToAXI4_xor281 ^ TLToAXI4_xor282;
  assign TLToAXI4_xor69 = TLToAXI4_xor139 ^ TLToAXI4_xor140;
  assign TLToAXI4_xor283 = count_64_pad ^ count_223_pad;
  assign TLToAXI4_xor284 = count_352_pad ^ count_153_pad;
  assign TLToAXI4_xor141 = TLToAXI4_xor283 ^ TLToAXI4_xor284;
  assign TLToAXI4_xor285 = count_118_pad ^ count_139_pad;
  assign TLToAXI4_xor286 = count_467_pad ^ count_386_pad;
  assign TLToAXI4_xor142 = TLToAXI4_xor285 ^ TLToAXI4_xor286;
  assign TLToAXI4_xor70 = TLToAXI4_xor141 ^ TLToAXI4_xor142;
  assign TLToAXI4_xor34 = TLToAXI4_xor69 ^ TLToAXI4_xor70;
  assign TLToAXI4_xor16 = TLToAXI4_xor33 ^ TLToAXI4_xor34;
  assign TLToAXI4_xor7 = TLToAXI4_xor15 ^ TLToAXI4_xor16;
  assign TLToAXI4_xor287 = count_434_pad ^ count_51_pad;
  assign TLToAXI4_xor288 = count_129_pad ^ count_378_pad;
  assign TLToAXI4_xor143 = TLToAXI4_xor287 ^ TLToAXI4_xor288;
  assign TLToAXI4_xor289 = count_186_pad ^ count_101_pad;
  assign TLToAXI4_xor290 = count_229_pad ^ count_280_pad;
  assign TLToAXI4_xor144 = TLToAXI4_xor289 ^ TLToAXI4_xor290;
  assign TLToAXI4_xor71 = TLToAXI4_xor143 ^ TLToAXI4_xor144;
  assign TLToAXI4_xor291 = count_403_pad ^ count_330_pad;
  assign TLToAXI4_xor292 = count_398_pad ^ count_307_pad;
  assign TLToAXI4_xor145 = TLToAXI4_xor291 ^ TLToAXI4_xor292;
  assign TLToAXI4_xor293 = count_216_pad ^ count_400_pad;
  assign TLToAXI4_xor294 = count_304_pad ^ count_131_pad;
  assign TLToAXI4_xor146 = TLToAXI4_xor293 ^ TLToAXI4_xor294;
  assign TLToAXI4_xor72 = TLToAXI4_xor145 ^ TLToAXI4_xor146;
  assign TLToAXI4_xor35 = TLToAXI4_xor71 ^ TLToAXI4_xor72;
  assign TLToAXI4_xor295 = count_282_pad ^ count_35_pad;
  assign TLToAXI4_xor296 = count_428_pad ^ count_16_pad;
  assign TLToAXI4_xor147 = TLToAXI4_xor295 ^ TLToAXI4_xor296;
  assign TLToAXI4_xor297 = count_355_pad ^ count_110_pad;
  assign TLToAXI4_xor298 = count_367_pad ^ count_427_pad;
  assign TLToAXI4_xor148 = TLToAXI4_xor297 ^ TLToAXI4_xor298;
  assign TLToAXI4_xor73 = TLToAXI4_xor147 ^ TLToAXI4_xor148;
  assign TLToAXI4_xor299 = count_46_pad ^ count_272_pad;
  assign TLToAXI4_xor300 = count_5_pad ^ count_173_pad;
  assign TLToAXI4_xor149 = TLToAXI4_xor299 ^ TLToAXI4_xor300;
  assign TLToAXI4_xor301 = count_211_pad ^ count_230_pad;
  assign TLToAXI4_xor302 = count_454_pad ^ count_458_pad;
  assign TLToAXI4_xor150 = TLToAXI4_xor301 ^ TLToAXI4_xor302;
  assign TLToAXI4_xor74 = TLToAXI4_xor149 ^ TLToAXI4_xor150;
  assign TLToAXI4_xor36 = TLToAXI4_xor73 ^ TLToAXI4_xor74;
  assign TLToAXI4_xor17 = TLToAXI4_xor35 ^ TLToAXI4_xor36;
  assign TLToAXI4_xor303 = count_23_pad ^ count_350_pad;
  assign TLToAXI4_xor304 = count_368_pad ^ count_456_pad;
  assign TLToAXI4_xor151 = TLToAXI4_xor303 ^ TLToAXI4_xor304;
  assign TLToAXI4_xor305 = count_464_pad ^ count_56_pad;
  assign TLToAXI4_xor306 = count_158_pad ^ count_1_pad;
  assign TLToAXI4_xor152 = TLToAXI4_xor305 ^ TLToAXI4_xor306;
  assign TLToAXI4_xor75 = TLToAXI4_xor151 ^ TLToAXI4_xor152;
  assign TLToAXI4_xor307 = count_62_pad ^ count_295_pad;
  assign TLToAXI4_xor308 = count_285_pad ^ count_44_pad;
  assign TLToAXI4_xor153 = TLToAXI4_xor307 ^ TLToAXI4_xor308;
  assign TLToAXI4_xor309 = count_25_pad ^ count_256_pad;
  assign TLToAXI4_xor310 = count_366_pad ^ count_473_pad;
  assign TLToAXI4_xor154 = TLToAXI4_xor309 ^ TLToAXI4_xor310;
  assign TLToAXI4_xor76 = TLToAXI4_xor153 ^ TLToAXI4_xor154;
  assign TLToAXI4_xor37 = TLToAXI4_xor75 ^ TLToAXI4_xor76;
  assign TLToAXI4_xor311 = count_465_pad ^ count_268_pad;
  assign TLToAXI4_xor312 = count_142_pad ^ count_75_pad;
  assign TLToAXI4_xor155 = TLToAXI4_xor311 ^ TLToAXI4_xor312;
  assign TLToAXI4_xor313 = count_240_pad ^ count_481_pad;
  assign TLToAXI4_xor314 = count_189_pad ^ count_382_pad;
  assign TLToAXI4_xor156 = TLToAXI4_xor313 ^ TLToAXI4_xor314;
  assign TLToAXI4_xor77 = TLToAXI4_xor155 ^ TLToAXI4_xor156;
  assign TLToAXI4_xor315 = count_219_pad ^ count_365_pad;
  assign TLToAXI4_xor316 = count_300_pad ^ count_53_pad;
  assign TLToAXI4_xor157 = TLToAXI4_xor315 ^ TLToAXI4_xor316;
  assign TLToAXI4_xor317 = count_490_pad ^ count_190_pad;
  assign TLToAXI4_xor638 = count_258_pad ^ count_356_pad;
  assign TLToAXI4_xor318 = count_332_pad ^ TLToAXI4_xor638;
  assign TLToAXI4_xor158 = TLToAXI4_xor317 ^ TLToAXI4_xor318;
  assign TLToAXI4_xor78 = TLToAXI4_xor157 ^ TLToAXI4_xor158;
  assign TLToAXI4_xor38 = TLToAXI4_xor77 ^ TLToAXI4_xor78;
  assign TLToAXI4_xor18 = TLToAXI4_xor37 ^ TLToAXI4_xor38;
  assign TLToAXI4_xor8 = TLToAXI4_xor17 ^ TLToAXI4_xor18;
  assign TLToAXI4_xor3 = TLToAXI4_xor7 ^ TLToAXI4_xor8;
  assign TLToAXI4_xor319 = count_410_pad ^ count_68_pad;
  assign TLToAXI4_xor320 = count_444_pad ^ count_446_pad;
  assign TLToAXI4_xor159 = TLToAXI4_xor319 ^ TLToAXI4_xor320;
  assign TLToAXI4_xor321 = count_493_pad ^ count_404_pad;
  assign TLToAXI4_xor322 = count_40_pad ^ count_495_pad;
  assign TLToAXI4_xor160 = TLToAXI4_xor321 ^ TLToAXI4_xor322;
  assign TLToAXI4_xor79 = TLToAXI4_xor159 ^ TLToAXI4_xor160;
  assign TLToAXI4_xor323 = count_325_pad ^ count_58_pad;
  assign TLToAXI4_xor324 = count_201_pad ^ count_107_pad;
  assign TLToAXI4_xor161 = TLToAXI4_xor323 ^ TLToAXI4_xor324;
  assign TLToAXI4_xor325 = count_292_pad ^ count_462_pad;
  assign TLToAXI4_xor326 = count_380_pad ^ count_57_pad;
  assign TLToAXI4_xor162 = TLToAXI4_xor325 ^ TLToAXI4_xor326;
  assign TLToAXI4_xor80 = TLToAXI4_xor161 ^ TLToAXI4_xor162;
  assign TLToAXI4_xor39 = TLToAXI4_xor79 ^ TLToAXI4_xor80;
  assign TLToAXI4_xor327 = count_395_pad ^ count_20_pad;
  assign TLToAXI4_xor328 = count_99_pad ^ count_327_pad;
  assign TLToAXI4_xor163 = TLToAXI4_xor327 ^ TLToAXI4_xor328;
  assign TLToAXI4_xor329 = count_30_pad ^ count_302_pad;
  assign TLToAXI4_xor330 = count_77_pad ^ count_439_pad;
  assign TLToAXI4_xor164 = TLToAXI4_xor329 ^ TLToAXI4_xor330;
  assign TLToAXI4_xor81 = TLToAXI4_xor163 ^ TLToAXI4_xor164;
  assign TLToAXI4_xor331 = count_409_pad ^ count_443_pad;
  assign TLToAXI4_xor332 = count_143_pad ^ count_165_pad;
  assign TLToAXI4_xor165 = TLToAXI4_xor331 ^ TLToAXI4_xor332;
  assign TLToAXI4_xor333 = count_81_pad ^ count_346_pad;
  assign TLToAXI4_xor334 = count_314_pad ^ count_196_pad;
  assign TLToAXI4_xor166 = TLToAXI4_xor333 ^ TLToAXI4_xor334;
  assign TLToAXI4_xor82 = TLToAXI4_xor165 ^ TLToAXI4_xor166;
  assign TLToAXI4_xor40 = TLToAXI4_xor81 ^ TLToAXI4_xor82;
  assign TLToAXI4_xor19 = TLToAXI4_xor39 ^ TLToAXI4_xor40;
  assign TLToAXI4_xor335 = count_262_pad ^ count_402_pad;
  assign TLToAXI4_xor336 = count_87_pad ^ count_29_pad;
  assign TLToAXI4_xor167 = TLToAXI4_xor335 ^ TLToAXI4_xor336;
  assign TLToAXI4_xor337 = count_126_pad ^ count_318_pad;
  assign TLToAXI4_xor338 = count_66_pad ^ count_163_pad;
  assign TLToAXI4_xor168 = TLToAXI4_xor337 ^ TLToAXI4_xor338;
  assign TLToAXI4_xor83 = TLToAXI4_xor167 ^ TLToAXI4_xor168;
  assign TLToAXI4_xor339 = count_175_pad ^ count_71_pad;
  assign TLToAXI4_xor340 = count_80_pad ^ count_252_pad;
  assign TLToAXI4_xor169 = TLToAXI4_xor339 ^ TLToAXI4_xor340;
  assign TLToAXI4_xor341 = count_28_pad ^ count_502_pad;
  assign TLToAXI4_xor342 = count_459_pad ^ count_141_pad;
  assign TLToAXI4_xor170 = TLToAXI4_xor341 ^ TLToAXI4_xor342;
  assign TLToAXI4_xor84 = TLToAXI4_xor169 ^ TLToAXI4_xor170;
  assign TLToAXI4_xor41 = TLToAXI4_xor83 ^ TLToAXI4_xor84;
  assign TLToAXI4_xor343 = count_405_pad ^ count_511_pad;
  assign TLToAXI4_xor344 = count_254_pad ^ count_476_pad;
  assign TLToAXI4_xor171 = TLToAXI4_xor343 ^ TLToAXI4_xor344;
  assign TLToAXI4_xor345 = count_97_pad ^ count_448_pad;
  assign TLToAXI4_xor346 = count_193_pad ^ count_260_pad;
  assign TLToAXI4_xor172 = TLToAXI4_xor345 ^ TLToAXI4_xor346;
  assign TLToAXI4_xor85 = TLToAXI4_xor171 ^ TLToAXI4_xor172;
  assign TLToAXI4_xor347 = count_303_pad ^ count_177_pad;
  assign TLToAXI4_xor348 = count_470_pad ^ count_146_pad;
  assign TLToAXI4_xor173 = TLToAXI4_xor347 ^ TLToAXI4_xor348;
  assign TLToAXI4_xor349 = count_309_pad ^ count_213_pad;
  assign TLToAXI4_xor350 = count_343_pad ^ count_468_pad;
  assign TLToAXI4_xor174 = TLToAXI4_xor349 ^ TLToAXI4_xor350;
  assign TLToAXI4_xor86 = TLToAXI4_xor173 ^ TLToAXI4_xor174;
  assign TLToAXI4_xor42 = TLToAXI4_xor85 ^ TLToAXI4_xor86;
  assign TLToAXI4_xor20 = TLToAXI4_xor41 ^ TLToAXI4_xor42;
  assign TLToAXI4_xor9 = TLToAXI4_xor19 ^ TLToAXI4_xor20;
  assign TLToAXI4_xor351 = count_429_pad ^ count_244_pad;
  assign TLToAXI4_xor352 = count_69_pad ^ count_460_pad;
  assign TLToAXI4_xor175 = TLToAXI4_xor351 ^ TLToAXI4_xor352;
  assign TLToAXI4_xor353 = count_370_pad ^ count_125_pad;
  assign TLToAXI4_xor354 = count_290_pad ^ count_128_pad;
  assign TLToAXI4_xor176 = TLToAXI4_xor353 ^ TLToAXI4_xor354;
  assign TLToAXI4_xor87 = TLToAXI4_xor175 ^ TLToAXI4_xor176;
  assign TLToAXI4_xor355 = count_407_pad ^ count_198_pad;
  assign TLToAXI4_xor356 = count_140_pad ^ count_512_pad;
  assign TLToAXI4_xor177 = TLToAXI4_xor355 ^ TLToAXI4_xor356;
  assign TLToAXI4_xor357 = count_440_pad ^ count_362_pad;
  assign TLToAXI4_xor358 = count_480_pad ^ count_109_pad;
  assign TLToAXI4_xor178 = TLToAXI4_xor357 ^ TLToAXI4_xor358;
  assign TLToAXI4_xor88 = TLToAXI4_xor177 ^ TLToAXI4_xor178;
  assign TLToAXI4_xor43 = TLToAXI4_xor87 ^ TLToAXI4_xor88;
  assign TLToAXI4_xor359 = count_171_pad ^ count_414_pad;
  assign TLToAXI4_xor360 = count_267_pad ^ count_484_pad;
  assign TLToAXI4_xor179 = TLToAXI4_xor359 ^ TLToAXI4_xor360;
  assign TLToAXI4_xor361 = count_278_pad ^ count_39_pad;
  assign TLToAXI4_xor362 = count_360_pad ^ count_14_pad;
  assign TLToAXI4_xor180 = TLToAXI4_xor361 ^ TLToAXI4_xor362;
  assign TLToAXI4_xor89 = TLToAXI4_xor179 ^ TLToAXI4_xor180;
  assign TLToAXI4_xor363 = count_336_pad ^ count_108_pad;
  assign TLToAXI4_xor364 = count_45_pad ^ count_275_pad;
  assign TLToAXI4_xor181 = TLToAXI4_xor363 ^ TLToAXI4_xor364;
  assign TLToAXI4_xor365 = count_413_pad ^ count_52_pad;
  assign TLToAXI4_xor366 = count_41_pad ^ count_328_pad;
  assign TLToAXI4_xor182 = TLToAXI4_xor365 ^ TLToAXI4_xor366;
  assign TLToAXI4_xor90 = TLToAXI4_xor181 ^ TLToAXI4_xor182;
  assign TLToAXI4_xor44 = TLToAXI4_xor89 ^ TLToAXI4_xor90;
  assign TLToAXI4_xor21 = TLToAXI4_xor43 ^ TLToAXI4_xor44;
  assign TLToAXI4_xor367 = count_82_pad ^ count_4_pad;
  assign TLToAXI4_xor368 = count_299_pad ^ count_286_pad;
  assign TLToAXI4_xor183 = TLToAXI4_xor367 ^ TLToAXI4_xor368;
  assign TLToAXI4_xor369 = count_510_pad ^ count_96_pad;
  assign TLToAXI4_xor370 = count_203_pad ^ count_452_pad;
  assign TLToAXI4_xor184 = TLToAXI4_xor369 ^ TLToAXI4_xor370;
  assign TLToAXI4_xor91 = TLToAXI4_xor183 ^ TLToAXI4_xor184;
  assign TLToAXI4_xor371 = count_150_pad ^ count_385_pad;
  assign TLToAXI4_xor372 = count_156_pad ^ count_169_pad;
  assign TLToAXI4_xor185 = TLToAXI4_xor371 ^ TLToAXI4_xor372;
  assign TLToAXI4_xor373 = count_132_pad ^ count_225_pad;
  assign TLToAXI4_xor374 = count_341_pad ^ count_377_pad;
  assign TLToAXI4_xor186 = TLToAXI4_xor373 ^ TLToAXI4_xor374;
  assign TLToAXI4_xor92 = TLToAXI4_xor185 ^ TLToAXI4_xor186;
  assign TLToAXI4_xor45 = TLToAXI4_xor91 ^ TLToAXI4_xor92;
  assign TLToAXI4_xor375 = count_114_pad ^ count_294_pad;
  assign TLToAXI4_xor376 = count_79_pad ^ count_60_pad;
  assign TLToAXI4_xor187 = TLToAXI4_xor375 ^ TLToAXI4_xor376;
  assign TLToAXI4_xor377 = count_86_pad ^ count_399_pad;
  assign TLToAXI4_xor378 = count_279_pad ^ count_239_pad;
  assign TLToAXI4_xor188 = TLToAXI4_xor377 ^ TLToAXI4_xor378;
  assign TLToAXI4_xor93 = TLToAXI4_xor187 ^ TLToAXI4_xor188;
  assign TLToAXI4_xor379 = count_13_pad ^ count_337_pad;
  assign TLToAXI4_xor380 = count_19_pad ^ count_334_pad;
  assign TLToAXI4_xor189 = TLToAXI4_xor379 ^ TLToAXI4_xor380;
  assign TLToAXI4_xor381 = count_17_pad ^ count_72_pad;
  assign TLToAXI4_xor766 = count_419_pad ^ count_176_pad;
  assign TLToAXI4_xor382 = count_94_pad ^ TLToAXI4_xor766;
  assign TLToAXI4_xor190 = TLToAXI4_xor381 ^ TLToAXI4_xor382;
  assign TLToAXI4_xor94 = TLToAXI4_xor189 ^ TLToAXI4_xor190;
  assign TLToAXI4_xor46 = TLToAXI4_xor93 ^ TLToAXI4_xor94;
  assign TLToAXI4_xor22 = TLToAXI4_xor45 ^ TLToAXI4_xor46;
  assign TLToAXI4_xor10 = TLToAXI4_xor21 ^ TLToAXI4_xor22;
  assign TLToAXI4_xor4 = TLToAXI4_xor9 ^ TLToAXI4_xor10;
  assign TLToAXI4_xor1 = TLToAXI4_xor3 ^ TLToAXI4_xor4;
  assign TLToAXI4_xor383 = count_210_pad ^ count_78_pad;
  assign TLToAXI4_xor384 = count_104_pad ^ count_507_pad;
  assign TLToAXI4_xor191 = TLToAXI4_xor383 ^ TLToAXI4_xor384;
  assign TLToAXI4_xor385 = count_287_pad ^ count_208_pad;
  assign TLToAXI4_xor386 = count_345_pad ^ count_311_pad;
  assign TLToAXI4_xor192 = TLToAXI4_xor385 ^ TLToAXI4_xor386;
  assign TLToAXI4_xor95 = TLToAXI4_xor191 ^ TLToAXI4_xor192;
  assign TLToAXI4_xor387 = count_178_pad ^ count_89_pad;
  assign TLToAXI4_xor388 = count_266_pad ^ count_238_pad;
  assign TLToAXI4_xor193 = TLToAXI4_xor387 ^ TLToAXI4_xor388;
  assign TLToAXI4_xor389 = count_206_pad ^ count_103_pad;
  assign TLToAXI4_xor390 = count_85_pad ^ count_138_pad;
  assign TLToAXI4_xor194 = TLToAXI4_xor389 ^ TLToAXI4_xor390;
  assign TLToAXI4_xor96 = TLToAXI4_xor193 ^ TLToAXI4_xor194;
  assign TLToAXI4_xor47 = TLToAXI4_xor95 ^ TLToAXI4_xor96;
  assign TLToAXI4_xor391 = count_392_pad ^ count_271_pad;
  assign TLToAXI4_xor392 = count_445_pad ^ count_431_pad;
  assign TLToAXI4_xor195 = TLToAXI4_xor391 ^ TLToAXI4_xor392;
  assign TLToAXI4_xor393 = count_220_pad ^ count_160_pad;
  assign TLToAXI4_xor394 = count_183_pad ^ count_436_pad;
  assign TLToAXI4_xor196 = TLToAXI4_xor393 ^ TLToAXI4_xor394;
  assign TLToAXI4_xor97 = TLToAXI4_xor195 ^ TLToAXI4_xor196;
  assign TLToAXI4_xor395 = count_226_pad ^ count_136_pad;
  assign TLToAXI4_xor396 = count_42_pad ^ count_351_pad;
  assign TLToAXI4_xor197 = TLToAXI4_xor395 ^ TLToAXI4_xor396;
  assign TLToAXI4_xor397 = count_261_pad ^ count_221_pad;
  assign TLToAXI4_xor398 = count_152_pad ^ count_505_pad;
  assign TLToAXI4_xor198 = TLToAXI4_xor397 ^ TLToAXI4_xor398;
  assign TLToAXI4_xor98 = TLToAXI4_xor197 ^ TLToAXI4_xor198;
  assign TLToAXI4_xor48 = TLToAXI4_xor97 ^ TLToAXI4_xor98;
  assign TLToAXI4_xor23 = TLToAXI4_xor47 ^ TLToAXI4_xor48;
  assign TLToAXI4_xor399 = count_36_pad ^ count_232_pad;
  assign TLToAXI4_xor400 = count_479_pad ^ count_34_pad;
  assign TLToAXI4_xor199 = TLToAXI4_xor399 ^ TLToAXI4_xor400;
  assign TLToAXI4_xor401 = count_291_pad ^ count_246_pad;
  assign TLToAXI4_xor402 = count_9_pad ^ count_98_pad;
  assign TLToAXI4_xor200 = TLToAXI4_xor401 ^ TLToAXI4_xor402;
  assign TLToAXI4_xor99 = TLToAXI4_xor199 ^ TLToAXI4_xor200;
  assign TLToAXI4_xor403 = count_364_pad ^ count_451_pad;
  assign TLToAXI4_xor404 = count_426_pad ^ count_492_pad;
  assign TLToAXI4_xor201 = TLToAXI4_xor403 ^ TLToAXI4_xor404;
  assign TLToAXI4_xor405 = count_281_pad ^ count_494_pad;
  assign TLToAXI4_xor406 = count_340_pad ^ count_179_pad;
  assign TLToAXI4_xor202 = TLToAXI4_xor405 ^ TLToAXI4_xor406;
  assign TLToAXI4_xor100 = TLToAXI4_xor201 ^ TLToAXI4_xor202;
  assign TLToAXI4_xor49 = TLToAXI4_xor99 ^ TLToAXI4_xor100;
  assign TLToAXI4_xor407 = count_250_pad ^ count_249_pad;
  assign TLToAXI4_xor408 = count_59_pad ^ count_320_pad;
  assign TLToAXI4_xor203 = TLToAXI4_xor407 ^ TLToAXI4_xor408;
  assign TLToAXI4_xor409 = count_321_pad ^ count_449_pad;
  assign TLToAXI4_xor410 = count_2_pad ^ count_496_pad;
  assign TLToAXI4_xor204 = TLToAXI4_xor409 ^ TLToAXI4_xor410;
  assign TLToAXI4_xor101 = TLToAXI4_xor203 ^ TLToAXI4_xor204;
  assign TLToAXI4_xor411 = count_188_pad ^ count_466_pad;
  assign TLToAXI4_xor412 = count_212_pad ^ count_11_pad;
  assign TLToAXI4_xor205 = TLToAXI4_xor411 ^ TLToAXI4_xor412;
  assign TLToAXI4_xor413 = count_55_pad ^ count_119_pad;
  assign TLToAXI4_xor414 = count_149_pad ^ count_450_pad;
  assign TLToAXI4_xor206 = TLToAXI4_xor413 ^ TLToAXI4_xor414;
  assign TLToAXI4_xor102 = TLToAXI4_xor205 ^ TLToAXI4_xor206;
  assign TLToAXI4_xor50 = TLToAXI4_xor101 ^ TLToAXI4_xor102;
  assign TLToAXI4_xor24 = TLToAXI4_xor49 ^ TLToAXI4_xor50;
  assign TLToAXI4_xor11 = TLToAXI4_xor23 ^ TLToAXI4_xor24;
  assign TLToAXI4_xor415 = count_32_pad ^ count_319_pad;
  assign TLToAXI4_xor416 = count_384_pad ^ count_162_pad;
  assign TLToAXI4_xor207 = TLToAXI4_xor415 ^ TLToAXI4_xor416;
  assign TLToAXI4_xor417 = count_231_pad ^ count_63_pad;
  assign TLToAXI4_xor418 = count_489_pad ^ count_509_pad;
  assign TLToAXI4_xor208 = TLToAXI4_xor417 ^ TLToAXI4_xor418;
  assign TLToAXI4_xor103 = TLToAXI4_xor207 ^ TLToAXI4_xor208;
  assign TLToAXI4_xor419 = count_133_pad ^ count_415_pad;
  assign TLToAXI4_xor420 = count_323_pad ^ count_289_pad;
  assign TLToAXI4_xor209 = TLToAXI4_xor419 ^ TLToAXI4_xor420;
  assign TLToAXI4_xor421 = count_342_pad ^ count_408_pad;
  assign TLToAXI4_xor422 = count_22_pad ^ count_308_pad;
  assign TLToAXI4_xor210 = TLToAXI4_xor421 ^ TLToAXI4_xor422;
  assign TLToAXI4_xor104 = TLToAXI4_xor209 ^ TLToAXI4_xor210;
  assign TLToAXI4_xor51 = TLToAXI4_xor103 ^ TLToAXI4_xor104;
  assign TLToAXI4_xor423 = count_424_pad ^ count_353_pad;
  assign TLToAXI4_xor424 = count_217_pad ^ count_497_pad;
  assign TLToAXI4_xor211 = TLToAXI4_xor423 ^ TLToAXI4_xor424;
  assign TLToAXI4_xor425 = count_430_pad ^ count_369_pad;
  assign TLToAXI4_xor426 = count_463_pad ^ count_389_pad;
  assign TLToAXI4_xor212 = TLToAXI4_xor425 ^ TLToAXI4_xor426;
  assign TLToAXI4_xor105 = TLToAXI4_xor211 ^ TLToAXI4_xor212;
  assign TLToAXI4_xor427 = count_499_pad ^ count_315_pad;
  assign TLToAXI4_xor428 = count_113_pad ^ count_506_pad;
  assign TLToAXI4_xor213 = TLToAXI4_xor427 ^ TLToAXI4_xor428;
  assign TLToAXI4_xor429 = count_257_pad ^ count_12_pad;
  assign TLToAXI4_xor430 = count_397_pad ^ count_326_pad;
  assign TLToAXI4_xor214 = TLToAXI4_xor429 ^ TLToAXI4_xor430;
  assign TLToAXI4_xor106 = TLToAXI4_xor213 ^ TLToAXI4_xor214;
  assign TLToAXI4_xor52 = TLToAXI4_xor105 ^ TLToAXI4_xor106;
  assign TLToAXI4_xor25 = TLToAXI4_xor51 ^ TLToAXI4_xor52;
  assign TLToAXI4_xor431 = count_469_pad ^ count_316_pad;
  assign TLToAXI4_xor432 = count_248_pad ^ r_first_pad;
  assign TLToAXI4_xor215 = TLToAXI4_xor431 ^ TLToAXI4_xor432;
  assign TLToAXI4_xor433 = count_390_pad ^ count_277_pad;
  assign TLToAXI4_xor434 = count_269_pad ^ count_218_pad;
  assign TLToAXI4_xor216 = TLToAXI4_xor433 ^ TLToAXI4_xor434;
  assign TLToAXI4_xor107 = TLToAXI4_xor215 ^ TLToAXI4_xor216;
  assign TLToAXI4_xor435 = count_115_pad ^ count_166_pad;
  assign TLToAXI4_xor436 = count_487_pad ^ count_192_pad;
  assign TLToAXI4_xor217 = TLToAXI4_xor435 ^ TLToAXI4_xor436;
  assign TLToAXI4_xor437 = count_508_pad ^ count_358_pad;
  assign TLToAXI4_xor438 = count_416_pad ^ count_151_pad;
  assign TLToAXI4_xor218 = TLToAXI4_xor437 ^ TLToAXI4_xor438;
  assign TLToAXI4_xor108 = TLToAXI4_xor217 ^ TLToAXI4_xor218;
  assign TLToAXI4_xor53 = TLToAXI4_xor107 ^ TLToAXI4_xor108;
  assign TLToAXI4_xor439 = count_354_pad ^ count_21_pad;
  assign TLToAXI4_xor440 = r_holds_d_pad ^ count_339_pad;
  assign TLToAXI4_xor219 = TLToAXI4_xor439 ^ TLToAXI4_xor440;
  assign TLToAXI4_xor441 = count_111_pad ^ count_18_pad;
  assign TLToAXI4_xor442 = count_425_pad ^ count_455_pad;
  assign TLToAXI4_xor220 = TLToAXI4_xor441 ^ TLToAXI4_xor442;
  assign TLToAXI4_xor109 = TLToAXI4_xor219 ^ TLToAXI4_xor220;
  assign TLToAXI4_xor443 = count_437_pad ^ count_245_pad;
  assign TLToAXI4_xor444 = count_116_pad ^ count_194_pad;
  assign TLToAXI4_xor221 = TLToAXI4_xor443 ^ TLToAXI4_xor444;
  assign TLToAXI4_xor445 = count_127_pad ^ count_137_pad;
  assign TLToAXI4_xor894 = count_159_pad ^ count_301_pad;
  assign TLToAXI4_xor446 = count_483_pad ^ TLToAXI4_xor894;
  assign TLToAXI4_xor222 = TLToAXI4_xor445 ^ TLToAXI4_xor446;
  assign TLToAXI4_xor110 = TLToAXI4_xor221 ^ TLToAXI4_xor222;
  assign TLToAXI4_xor54 = TLToAXI4_xor109 ^ TLToAXI4_xor110;
  assign TLToAXI4_xor26 = TLToAXI4_xor53 ^ TLToAXI4_xor54;
  assign TLToAXI4_xor12 = TLToAXI4_xor25 ^ TLToAXI4_xor26;
  assign TLToAXI4_xor5 = TLToAXI4_xor11 ^ TLToAXI4_xor12;
  assign TLToAXI4_xor447 = count_215_pad ^ count_288_pad;
  assign TLToAXI4_xor448 = count_54_pad ^ count_27_pad;
  assign TLToAXI4_xor223 = TLToAXI4_xor447 ^ TLToAXI4_xor448;
  assign TLToAXI4_xor449 = count_161_pad ^ count_106_pad;
  assign TLToAXI4_xor450 = count_485_pad ^ count_259_pad;
  assign TLToAXI4_xor224 = TLToAXI4_xor449 ^ TLToAXI4_xor450;
  assign TLToAXI4_xor111 = TLToAXI4_xor223 ^ TLToAXI4_xor224;
  assign TLToAXI4_xor451 = count_264_pad ^ count_91_pad;
  assign TLToAXI4_xor452 = count_84_pad ^ count_312_pad;
  assign TLToAXI4_xor225 = TLToAXI4_xor451 ^ TLToAXI4_xor452;
  assign TLToAXI4_xor453 = count_207_pad ^ count_172_pad;
  assign TLToAXI4_xor454 = count_253_pad ^ count_148_pad;
  assign TLToAXI4_xor226 = TLToAXI4_xor453 ^ TLToAXI4_xor454;
  assign TLToAXI4_xor112 = TLToAXI4_xor225 ^ TLToAXI4_xor226;
  assign TLToAXI4_xor55 = TLToAXI4_xor111 ^ TLToAXI4_xor112;
  assign TLToAXI4_xor455 = count_228_pad ^ count_10_pad;
  assign TLToAXI4_xor456 = count_322_pad ^ count_363_pad;
  assign TLToAXI4_xor227 = TLToAXI4_xor455 ^ TLToAXI4_xor456;
  assign TLToAXI4_xor457 = count_48_pad ^ count_236_pad;
  assign TLToAXI4_xor458 = count_205_pad ^ count_191_pad;
  assign TLToAXI4_xor228 = TLToAXI4_xor457 ^ TLToAXI4_xor458;
  assign TLToAXI4_xor113 = TLToAXI4_xor227 ^ TLToAXI4_xor228;
  assign TLToAXI4_xor459 = count_338_pad ^ count_276_pad;
  assign TLToAXI4_xor460 = count_475_pad ^ count_24_pad;
  assign TLToAXI4_xor229 = TLToAXI4_xor459 ^ TLToAXI4_xor460;
  assign TLToAXI4_xor461 = count_387_pad ^ count_438_pad;
  assign TLToAXI4_xor462 = count_472_pad ^ count_167_pad;
  assign TLToAXI4_xor230 = TLToAXI4_xor461 ^ TLToAXI4_xor462;
  assign TLToAXI4_xor114 = TLToAXI4_xor229 ^ TLToAXI4_xor230;
  assign TLToAXI4_xor56 = TLToAXI4_xor113 ^ TLToAXI4_xor114;
  assign TLToAXI4_xor27 = TLToAXI4_xor55 ^ TLToAXI4_xor56;
  assign TLToAXI4_xor463 = count_233_pad ^ count_185_pad;
  assign TLToAXI4_xor464 = count_135_pad ^ count_197_pad;
  assign TLToAXI4_xor231 = TLToAXI4_xor463 ^ TLToAXI4_xor464;
  assign TLToAXI4_xor465 = count_273_pad ^ count_441_pad;
  assign TLToAXI4_xor466 = count_88_pad ^ count_471_pad;
  assign TLToAXI4_xor232 = TLToAXI4_xor465 ^ TLToAXI4_xor466;
  assign TLToAXI4_xor115 = TLToAXI4_xor231 ^ TLToAXI4_xor232;
  assign TLToAXI4_xor467 = count_147_pad ^ count_412_pad;
  assign TLToAXI4_xor468 = count_488_pad ^ count_486_pad;
  assign TLToAXI4_xor233 = TLToAXI4_xor467 ^ TLToAXI4_xor468;
  assign TLToAXI4_xor469 = count_298_pad ^ count_442_pad;
  assign TLToAXI4_xor470 = count_73_pad ^ count_237_pad;
  assign TLToAXI4_xor234 = TLToAXI4_xor469 ^ TLToAXI4_xor470;
  assign TLToAXI4_xor116 = TLToAXI4_xor233 ^ TLToAXI4_xor234;
  assign TLToAXI4_xor57 = TLToAXI4_xor115 ^ TLToAXI4_xor116;
  assign TLToAXI4_xor471 = count_435_pad ^ count_6_pad;
  assign TLToAXI4_xor472 = count_361_pad ^ count_15_pad;
  assign TLToAXI4_xor235 = TLToAXI4_xor471 ^ TLToAXI4_xor472;
  assign TLToAXI4_xor473 = count_388_pad ^ count_164_pad;
  assign TLToAXI4_xor474 = count_255_pad ^ count_306_pad;
  assign TLToAXI4_xor236 = TLToAXI4_xor473 ^ TLToAXI4_xor474;
  assign TLToAXI4_xor117 = TLToAXI4_xor235 ^ TLToAXI4_xor236;
  assign TLToAXI4_xor475 = count_381_pad ^ count_130_pad;
  assign TLToAXI4_xor476 = count_145_pad ^ count_8_pad;
  assign TLToAXI4_xor237 = TLToAXI4_xor475 ^ TLToAXI4_xor476;
  assign TLToAXI4_xor477 = count_224_pad ^ count_349_pad;
  assign TLToAXI4_xor478 = count_375_pad ^ count_457_pad;
  assign TLToAXI4_xor238 = TLToAXI4_xor477 ^ TLToAXI4_xor478;
  assign TLToAXI4_xor118 = TLToAXI4_xor237 ^ TLToAXI4_xor238;
  assign TLToAXI4_xor58 = TLToAXI4_xor117 ^ TLToAXI4_xor118;
  assign TLToAXI4_xor28 = TLToAXI4_xor57 ^ TLToAXI4_xor58;
  assign TLToAXI4_xor13 = TLToAXI4_xor27 ^ TLToAXI4_xor28;
  assign TLToAXI4_xor479 = b_delay_pad ^ count_181_pad;
  assign TLToAXI4_xor480 = count_170_pad ^ count_3_pad;
  assign TLToAXI4_xor239 = TLToAXI4_xor479 ^ TLToAXI4_xor480;
  assign TLToAXI4_xor481 = count_461_pad ^ count_102_pad;
  assign TLToAXI4_xor482 = count_134_pad ^ count_234_pad;
  assign TLToAXI4_xor240 = TLToAXI4_xor481 ^ TLToAXI4_xor482;
  assign TLToAXI4_xor119 = TLToAXI4_xor239 ^ TLToAXI4_xor240;
  assign TLToAXI4_xor483 = count_335_pad ^ count_95_pad;
  assign TLToAXI4_xor484 = count_374_pad ^ count_49_pad;
  assign TLToAXI4_xor241 = TLToAXI4_xor483 ^ TLToAXI4_xor484;
  assign TLToAXI4_xor485 = count_100_pad ^ count_283_pad;
  assign TLToAXI4_xor486 = count_90_pad ^ count_155_pad;
  assign TLToAXI4_xor242 = TLToAXI4_xor485 ^ TLToAXI4_xor486;
  assign TLToAXI4_xor120 = TLToAXI4_xor241 ^ TLToAXI4_xor242;
  assign TLToAXI4_xor59 = TLToAXI4_xor119 ^ TLToAXI4_xor120;
  assign TLToAXI4_xor487 = count_274_pad ^ count_83_pad;
  assign TLToAXI4_xor488 = count_112_pad ^ count_433_pad;
  assign TLToAXI4_xor243 = TLToAXI4_xor487 ^ TLToAXI4_xor488;
  assign TLToAXI4_xor489 = count_93_pad ^ count_65_pad;
  assign TLToAXI4_xor490 = count_235_pad ^ count_371_pad;
  assign TLToAXI4_xor244 = TLToAXI4_xor489 ^ TLToAXI4_xor490;
  assign TLToAXI4_xor121 = TLToAXI4_xor243 ^ TLToAXI4_xor244;
  assign TLToAXI4_xor491 = count_122_pad ^ count_247_pad;
  assign TLToAXI4_xor492 = count_157_pad ^ count_180_pad;
  assign TLToAXI4_xor245 = TLToAXI4_xor491 ^ TLToAXI4_xor492;
  assign TLToAXI4_xor493 = count_347_pad ^ count_251_pad;
  assign TLToAXI4_xor494 = count_200_pad ^ count_187_pad;
  assign TLToAXI4_xor246 = TLToAXI4_xor493 ^ TLToAXI4_xor494;
  assign TLToAXI4_xor122 = TLToAXI4_xor245 ^ TLToAXI4_xor246;
  assign TLToAXI4_xor60 = TLToAXI4_xor121 ^ TLToAXI4_xor122;
  assign TLToAXI4_xor29 = TLToAXI4_xor59 ^ TLToAXI4_xor60;
  assign TLToAXI4_xor495 = count_432_pad ^ count_123_pad;
  assign TLToAXI4_xor496 = count_418_pad ^ count_406_pad;
  assign TLToAXI4_xor247 = TLToAXI4_xor495 ^ TLToAXI4_xor496;
  assign TLToAXI4_xor497 = count_241_pad ^ count_33_pad;
  assign TLToAXI4_xor498 = count_324_pad ^ count_105_pad;
  assign TLToAXI4_xor248 = TLToAXI4_xor497 ^ TLToAXI4_xor498;
  assign TLToAXI4_xor123 = TLToAXI4_xor247 ^ TLToAXI4_xor248;
  assign TLToAXI4_xor499 = count_92_pad ^ count_7_pad;
  assign TLToAXI4_xor500 = count_214_pad ^ count_379_pad;
  assign TLToAXI4_xor249 = TLToAXI4_xor499 ^ TLToAXI4_xor500;
  assign TLToAXI4_xor501 = count_359_pad ^ doneAW_pad;
  assign TLToAXI4_xor502 = count_144_pad ^ count_396_pad;
  assign TLToAXI4_xor250 = TLToAXI4_xor501 ^ TLToAXI4_xor502;
  assign TLToAXI4_xor124 = TLToAXI4_xor249 ^ TLToAXI4_xor250;
  assign TLToAXI4_xor61 = TLToAXI4_xor123 ^ TLToAXI4_xor124;
  assign TLToAXI4_xor503 = count_376_pad ^ count_504_pad;
  assign TLToAXI4_xor504 = count_124_pad ^ count_500_pad;
  assign TLToAXI4_xor251 = TLToAXI4_xor503 ^ TLToAXI4_xor504;
  assign TLToAXI4_xor505 = count_209_pad ^ count_348_pad;
  assign TLToAXI4_xor506 = count_344_pad ^ count_76_pad;
  assign TLToAXI4_xor252 = TLToAXI4_xor505 ^ TLToAXI4_xor506;
  assign TLToAXI4_xor125 = TLToAXI4_xor251 ^ TLToAXI4_xor252;
  assign TLToAXI4_xor507 = count_265_pad ^ count_453_pad;
  assign TLToAXI4_xor508 = count_47_pad ^ count_43_pad;
  assign TLToAXI4_xor253 = TLToAXI4_xor507 ^ TLToAXI4_xor508;
  assign TLToAXI4_xor509 = count_74_pad ^ count_491_pad;
  assign TLToAXI4_xor1022 = count_243_pad ^ count_174_pad;
  assign TLToAXI4_xor510 = count_478_pad ^ TLToAXI4_xor1022;
  assign TLToAXI4_xor254 = TLToAXI4_xor509 ^ TLToAXI4_xor510;
  assign TLToAXI4_xor126 = TLToAXI4_xor253 ^ TLToAXI4_xor254;
  assign TLToAXI4_xor62 = TLToAXI4_xor125 ^ TLToAXI4_xor126;
  assign TLToAXI4_xor30 = TLToAXI4_xor61 ^ TLToAXI4_xor62;
  assign TLToAXI4_xor14 = TLToAXI4_xor29 ^ TLToAXI4_xor30;
  assign TLToAXI4_xor6 = TLToAXI4_xor13 ^ TLToAXI4_xor14;
  assign TLToAXI4_xor2 = TLToAXI4_xor5 ^ TLToAXI4_xor6;
  assign TLToAXI4_xor0 = TLToAXI4_xor1 ^ TLToAXI4_xor2;
  assign deq_sum = TLToAXI4_covSum + deq_io_covSum;
  assign queue_arw_deq_sum = deq_sum + queue_arw_deq_io_covSum;
  assign io_covSum = queue_arw_deq_sum;
  assign deq_metaReset = metaReset;
  assign queue_arw_deq_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_512 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_512 <= count_512 + inc_511 - dec_511; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_511 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_511 <= count_511 + inc_510 - dec_510; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_510 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_510 <= count_510 + inc_509 - dec_509; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_509 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_509 <= count_509 + inc_508 - dec_508; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_508 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_508 <= count_508 + inc_507 - dec_507; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_507 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_507 <= count_507 + inc_506 - dec_506; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_506 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_506 <= count_506 + inc_505 - dec_505; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_505 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_505 <= count_505 + inc_504 - dec_504; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_504 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_504 <= count_504 + inc_503 - dec_503; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_503 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_503 <= count_503 + inc_502 - dec_502; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_502 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_502 <= count_502 + inc_501 - dec_501; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_501 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_501 <= count_501 + inc_500 - dec_500; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_500 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_500 <= count_500 + inc_499 - dec_499; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_499 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_499 <= count_499 + inc_498 - dec_498; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_498 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_498 <= count_498 + inc_497 - dec_497; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_497 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_497 <= count_497 + inc_496 - dec_496; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_496 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_496 <= count_496 + inc_495 - dec_495; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_495 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_495 <= count_495 + inc_494 - dec_494; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_494 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_494 <= count_494 + inc_493 - dec_493; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_493 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_493 <= count_493 + inc_492 - dec_492; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_492 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_492 <= count_492 + inc_491 - dec_491; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_491 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_491 <= count_491 + inc_490 - dec_490; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_490 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_490 <= count_490 + inc_489 - dec_489; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_489 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_489 <= count_489 + inc_488 - dec_488; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_488 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_488 <= count_488 + inc_487 - dec_487; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_487 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_487 <= count_487 + inc_486 - dec_486; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_486 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_486 <= count_486 + inc_485 - dec_485; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_485 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_485 <= count_485 + inc_484 - dec_484; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_484 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_484 <= count_484 + inc_483 - dec_483; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_483 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_483 <= count_483 + inc_482 - dec_482; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_482 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_482 <= count_482 + inc_481 - dec_481; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_481 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_481 <= count_481 + inc_480 - dec_480; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_480 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_480 <= count_480 + inc_479 - dec_479; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_479 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_479 <= count_479 + inc_478 - dec_478; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_478 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_478 <= count_478 + inc_477 - dec_477; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_477 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_477 <= count_477 + inc_476 - dec_476; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_476 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_476 <= count_476 + inc_475 - dec_475; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_475 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_475 <= count_475 + inc_474 - dec_474; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_474 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_474 <= count_474 + inc_473 - dec_473; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_473 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_473 <= count_473 + inc_472 - dec_472; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_472 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_472 <= count_472 + inc_471 - dec_471; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_471 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_471 <= count_471 + inc_470 - dec_470; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_470 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_470 <= count_470 + inc_469 - dec_469; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_469 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_469 <= count_469 + inc_468 - dec_468; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_468 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_468 <= count_468 + inc_467 - dec_467; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_467 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_467 <= count_467 + inc_466 - dec_466; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_466 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_466 <= count_466 + inc_465 - dec_465; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_465 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_465 <= count_465 + inc_464 - dec_464; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_464 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_464 <= count_464 + inc_463 - dec_463; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_463 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_463 <= count_463 + inc_462 - dec_462; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_462 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_462 <= count_462 + inc_461 - dec_461; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_461 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_461 <= count_461 + inc_460 - dec_460; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_460 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_460 <= count_460 + inc_459 - dec_459; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_459 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_459 <= count_459 + inc_458 - dec_458; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_458 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_458 <= count_458 + inc_457 - dec_457; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_457 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_457 <= count_457 + inc_456 - dec_456; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_456 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_456 <= count_456 + inc_455 - dec_455; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_455 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_455 <= count_455 + inc_454 - dec_454; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_454 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_454 <= count_454 + inc_453 - dec_453; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_453 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_453 <= count_453 + inc_452 - dec_452; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_452 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_452 <= count_452 + inc_451 - dec_451; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_451 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_451 <= count_451 + inc_450 - dec_450; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_450 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_450 <= count_450 + inc_449 - dec_449; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_449 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_449 <= count_449 + inc_448 - dec_448; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_448 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_448 <= count_448 + inc_447 - dec_447; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_447 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_447 <= count_447 + inc_446 - dec_446; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_446 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_446 <= count_446 + inc_445 - dec_445; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_445 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_445 <= count_445 + inc_444 - dec_444; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_444 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_444 <= count_444 + inc_443 - dec_443; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_443 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_443 <= count_443 + inc_442 - dec_442; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_442 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_442 <= count_442 + inc_441 - dec_441; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_441 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_441 <= count_441 + inc_440 - dec_440; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_440 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_440 <= count_440 + inc_439 - dec_439; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_439 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_439 <= count_439 + inc_438 - dec_438; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_438 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_438 <= count_438 + inc_437 - dec_437; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_437 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_437 <= count_437 + inc_436 - dec_436; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_436 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_436 <= count_436 + inc_435 - dec_435; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_435 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_435 <= count_435 + inc_434 - dec_434; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_434 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_434 <= count_434 + inc_433 - dec_433; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_433 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_433 <= count_433 + inc_432 - dec_432; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_432 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_432 <= count_432 + inc_431 - dec_431; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_431 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_431 <= count_431 + inc_430 - dec_430; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_430 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_430 <= count_430 + inc_429 - dec_429; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_429 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_429 <= count_429 + inc_428 - dec_428; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_428 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_428 <= count_428 + inc_427 - dec_427; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_427 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_427 <= count_427 + inc_426 - dec_426; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_426 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_426 <= count_426 + inc_425 - dec_425; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_425 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_425 <= count_425 + inc_424 - dec_424; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_424 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_424 <= count_424 + inc_423 - dec_423; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_423 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_423 <= count_423 + inc_422 - dec_422; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_422 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_422 <= count_422 + inc_421 - dec_421; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_421 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_421 <= count_421 + inc_420 - dec_420; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_420 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_420 <= count_420 + inc_419 - dec_419; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_419 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_419 <= count_419 + inc_418 - dec_418; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_418 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_418 <= count_418 + inc_417 - dec_417; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_417 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_417 <= count_417 + inc_416 - dec_416; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_416 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_416 <= count_416 + inc_415 - dec_415; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_415 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_415 <= count_415 + inc_414 - dec_414; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_414 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_414 <= count_414 + inc_413 - dec_413; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_413 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_413 <= count_413 + inc_412 - dec_412; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_412 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_412 <= count_412 + inc_411 - dec_411; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_411 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_411 <= count_411 + inc_410 - dec_410; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_410 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_410 <= count_410 + inc_409 - dec_409; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_409 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_409 <= count_409 + inc_408 - dec_408; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_408 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_408 <= count_408 + inc_407 - dec_407; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_407 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_407 <= count_407 + inc_406 - dec_406; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_406 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_406 <= count_406 + inc_405 - dec_405; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_405 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_405 <= count_405 + inc_404 - dec_404; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_404 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_404 <= count_404 + inc_403 - dec_403; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_403 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_403 <= count_403 + inc_402 - dec_402; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_402 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_402 <= count_402 + inc_401 - dec_401; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_401 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_401 <= count_401 + inc_400 - dec_400; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_400 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_400 <= count_400 + inc_399 - dec_399; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_399 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_399 <= count_399 + inc_398 - dec_398; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_398 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_398 <= count_398 + inc_397 - dec_397; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_397 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_397 <= count_397 + inc_396 - dec_396; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_396 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_396 <= count_396 + inc_395 - dec_395; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_395 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_395 <= count_395 + inc_394 - dec_394; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_394 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_394 <= count_394 + inc_393 - dec_393; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_393 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_393 <= count_393 + inc_392 - dec_392; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_392 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_392 <= count_392 + inc_391 - dec_391; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_391 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_391 <= count_391 + inc_390 - dec_390; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_390 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_390 <= count_390 + inc_389 - dec_389; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_389 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_389 <= count_389 + inc_388 - dec_388; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_388 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_388 <= count_388 + inc_387 - dec_387; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_387 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_387 <= count_387 + inc_386 - dec_386; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_386 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_386 <= count_386 + inc_385 - dec_385; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_385 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_385 <= count_385 + inc_384 - dec_384; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_384 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_384 <= count_384 + inc_383 - dec_383; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_383 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_383 <= count_383 + inc_382 - dec_382; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_382 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_382 <= count_382 + inc_381 - dec_381; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_381 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_381 <= count_381 + inc_380 - dec_380; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_380 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_380 <= count_380 + inc_379 - dec_379; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_379 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_379 <= count_379 + inc_378 - dec_378; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_378 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_378 <= count_378 + inc_377 - dec_377; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_377 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_377 <= count_377 + inc_376 - dec_376; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_376 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_376 <= count_376 + inc_375 - dec_375; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_375 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_375 <= count_375 + inc_374 - dec_374; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_374 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_374 <= count_374 + inc_373 - dec_373; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_373 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_373 <= count_373 + inc_372 - dec_372; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_372 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_372 <= count_372 + inc_371 - dec_371; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_371 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_371 <= count_371 + inc_370 - dec_370; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_370 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_370 <= count_370 + inc_369 - dec_369; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_369 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_369 <= count_369 + inc_368 - dec_368; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_368 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_368 <= count_368 + inc_367 - dec_367; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_367 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_367 <= count_367 + inc_366 - dec_366; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_366 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_366 <= count_366 + inc_365 - dec_365; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_365 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_365 <= count_365 + inc_364 - dec_364; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_364 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_364 <= count_364 + inc_363 - dec_363; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_363 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_363 <= count_363 + inc_362 - dec_362; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_362 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_362 <= count_362 + inc_361 - dec_361; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_361 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_361 <= count_361 + inc_360 - dec_360; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_360 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_360 <= count_360 + inc_359 - dec_359; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_359 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_359 <= count_359 + inc_358 - dec_358; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_358 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_358 <= count_358 + inc_357 - dec_357; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_357 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_357 <= count_357 + inc_356 - dec_356; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_356 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_356 <= count_356 + inc_355 - dec_355; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_355 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_355 <= count_355 + inc_354 - dec_354; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_354 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_354 <= count_354 + inc_353 - dec_353; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_353 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_353 <= count_353 + inc_352 - dec_352; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_352 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_352 <= count_352 + inc_351 - dec_351; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_351 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_351 <= count_351 + inc_350 - dec_350; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_350 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_350 <= count_350 + inc_349 - dec_349; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_349 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_349 <= count_349 + inc_348 - dec_348; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_348 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_348 <= count_348 + inc_347 - dec_347; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_347 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_347 <= count_347 + inc_346 - dec_346; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_346 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_346 <= count_346 + inc_345 - dec_345; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_345 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_345 <= count_345 + inc_344 - dec_344; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_344 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_344 <= count_344 + inc_343 - dec_343; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_343 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_343 <= count_343 + inc_342 - dec_342; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_342 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_342 <= count_342 + inc_341 - dec_341; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_341 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_341 <= count_341 + inc_340 - dec_340; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_340 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_340 <= count_340 + inc_339 - dec_339; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_339 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_339 <= count_339 + inc_338 - dec_338; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_338 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_338 <= count_338 + inc_337 - dec_337; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_337 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_337 <= count_337 + inc_336 - dec_336; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_336 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_336 <= count_336 + inc_335 - dec_335; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_335 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_335 <= count_335 + inc_334 - dec_334; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_334 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_334 <= count_334 + inc_333 - dec_333; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_333 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_333 <= count_333 + inc_332 - dec_332; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_332 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_332 <= count_332 + inc_331 - dec_331; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_331 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_331 <= count_331 + inc_330 - dec_330; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_330 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_330 <= count_330 + inc_329 - dec_329; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_329 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_329 <= count_329 + inc_328 - dec_328; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_328 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_328 <= count_328 + inc_327 - dec_327; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_327 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_327 <= count_327 + inc_326 - dec_326; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_326 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_326 <= count_326 + inc_325 - dec_325; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_325 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_325 <= count_325 + inc_324 - dec_324; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_324 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_324 <= count_324 + inc_323 - dec_323; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_323 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_323 <= count_323 + inc_322 - dec_322; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_322 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_322 <= count_322 + inc_321 - dec_321; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_321 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_321 <= count_321 + inc_320 - dec_320; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_320 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_320 <= count_320 + inc_319 - dec_319; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_319 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_319 <= count_319 + inc_318 - dec_318; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_318 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_318 <= count_318 + inc_317 - dec_317; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_317 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_317 <= count_317 + inc_316 - dec_316; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_316 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_316 <= count_316 + inc_315 - dec_315; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_315 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_315 <= count_315 + inc_314 - dec_314; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_314 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_314 <= count_314 + inc_313 - dec_313; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_313 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_313 <= count_313 + inc_312 - dec_312; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_312 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_312 <= count_312 + inc_311 - dec_311; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_311 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_311 <= count_311 + inc_310 - dec_310; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_310 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_310 <= count_310 + inc_309 - dec_309; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_309 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_309 <= count_309 + inc_308 - dec_308; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_308 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_308 <= count_308 + inc_307 - dec_307; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_307 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_307 <= count_307 + inc_306 - dec_306; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_306 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_306 <= count_306 + inc_305 - dec_305; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_305 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_305 <= count_305 + inc_304 - dec_304; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_304 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_304 <= count_304 + inc_303 - dec_303; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_303 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_303 <= count_303 + inc_302 - dec_302; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_302 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_302 <= count_302 + inc_301 - dec_301; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_301 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_301 <= count_301 + inc_300 - dec_300; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_300 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_300 <= count_300 + inc_299 - dec_299; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_299 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_299 <= count_299 + inc_298 - dec_298; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_298 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_298 <= count_298 + inc_297 - dec_297; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_297 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_297 <= count_297 + inc_296 - dec_296; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_296 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_296 <= count_296 + inc_295 - dec_295; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_295 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_295 <= count_295 + inc_294 - dec_294; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_294 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_294 <= count_294 + inc_293 - dec_293; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_293 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_293 <= count_293 + inc_292 - dec_292; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_292 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_292 <= count_292 + inc_291 - dec_291; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_291 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_291 <= count_291 + inc_290 - dec_290; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_290 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_290 <= count_290 + inc_289 - dec_289; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_289 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_289 <= count_289 + inc_288 - dec_288; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_288 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_288 <= count_288 + inc_287 - dec_287; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_287 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_287 <= count_287 + inc_286 - dec_286; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_286 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_286 <= count_286 + inc_285 - dec_285; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_285 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_285 <= count_285 + inc_284 - dec_284; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_284 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_284 <= count_284 + inc_283 - dec_283; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_283 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_283 <= count_283 + inc_282 - dec_282; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_282 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_282 <= count_282 + inc_281 - dec_281; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_281 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_281 <= count_281 + inc_280 - dec_280; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_280 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_280 <= count_280 + inc_279 - dec_279; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_279 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_279 <= count_279 + inc_278 - dec_278; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_278 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_278 <= count_278 + inc_277 - dec_277; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_277 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_277 <= count_277 + inc_276 - dec_276; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_276 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_276 <= count_276 + inc_275 - dec_275; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_275 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_275 <= count_275 + inc_274 - dec_274; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_274 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_274 <= count_274 + inc_273 - dec_273; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_273 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_273 <= count_273 + inc_272 - dec_272; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_272 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_272 <= count_272 + inc_271 - dec_271; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_271 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_271 <= count_271 + inc_270 - dec_270; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_270 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_270 <= count_270 + inc_269 - dec_269; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_269 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_269 <= count_269 + inc_268 - dec_268; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_268 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_268 <= count_268 + inc_267 - dec_267; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_267 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_267 <= count_267 + inc_266 - dec_266; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_266 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_266 <= count_266 + inc_265 - dec_265; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_265 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_265 <= count_265 + inc_264 - dec_264; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_264 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_264 <= count_264 + inc_263 - dec_263; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_263 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_263 <= count_263 + inc_262 - dec_262; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_262 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_262 <= count_262 + inc_261 - dec_261; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_261 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_261 <= count_261 + inc_260 - dec_260; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_260 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_260 <= count_260 + inc_259 - dec_259; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_259 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_259 <= count_259 + inc_258 - dec_258; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_258 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_258 <= count_258 + inc_257 - dec_257; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_257 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_257 <= count_257 + inc_256 - dec_256; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_256 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_256 <= count_256 + inc_255 - dec_255; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_255 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_255 <= count_255 + inc_254 - dec_254; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_254 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_254 <= count_254 + inc_253 - dec_253; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_253 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_253 <= count_253 + inc_252 - dec_252; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_252 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_252 <= count_252 + inc_251 - dec_251; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_251 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_251 <= count_251 + inc_250 - dec_250; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_250 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_250 <= count_250 + inc_249 - dec_249; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_249 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_249 <= count_249 + inc_248 - dec_248; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_248 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_248 <= count_248 + inc_247 - dec_247; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_247 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_247 <= count_247 + inc_246 - dec_246; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_246 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_246 <= count_246 + inc_245 - dec_245; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_245 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_245 <= count_245 + inc_244 - dec_244; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_244 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_244 <= count_244 + inc_243 - dec_243; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_243 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_243 <= count_243 + inc_242 - dec_242; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_242 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_242 <= count_242 + inc_241 - dec_241; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_241 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_241 <= count_241 + inc_240 - dec_240; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_240 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_240 <= count_240 + inc_239 - dec_239; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_239 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_239 <= count_239 + inc_238 - dec_238; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_238 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_238 <= count_238 + inc_237 - dec_237; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_237 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_237 <= count_237 + inc_236 - dec_236; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_236 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_236 <= count_236 + inc_235 - dec_235; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_235 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_235 <= count_235 + inc_234 - dec_234; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_234 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_234 <= count_234 + inc_233 - dec_233; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_233 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_233 <= count_233 + inc_232 - dec_232; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_232 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_232 <= count_232 + inc_231 - dec_231; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_231 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_231 <= count_231 + inc_230 - dec_230; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_230 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_230 <= count_230 + inc_229 - dec_229; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_229 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_229 <= count_229 + inc_228 - dec_228; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_228 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_228 <= count_228 + inc_227 - dec_227; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_227 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_227 <= count_227 + inc_226 - dec_226; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_226 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_226 <= count_226 + inc_225 - dec_225; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_225 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_225 <= count_225 + inc_224 - dec_224; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_224 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_224 <= count_224 + inc_223 - dec_223; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_223 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_223 <= count_223 + inc_222 - dec_222; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_222 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_222 <= count_222 + inc_221 - dec_221; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_221 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_221 <= count_221 + inc_220 - dec_220; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_220 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_220 <= count_220 + inc_219 - dec_219; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_219 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_219 <= count_219 + inc_218 - dec_218; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_218 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_218 <= count_218 + inc_217 - dec_217; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_217 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_217 <= count_217 + inc_216 - dec_216; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_216 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_216 <= count_216 + inc_215 - dec_215; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_215 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_215 <= count_215 + inc_214 - dec_214; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_214 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_214 <= count_214 + inc_213 - dec_213; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_213 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_213 <= count_213 + inc_212 - dec_212; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_212 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_212 <= count_212 + inc_211 - dec_211; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_211 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_211 <= count_211 + inc_210 - dec_210; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_210 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_210 <= count_210 + inc_209 - dec_209; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_209 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_209 <= count_209 + inc_208 - dec_208; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_208 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_208 <= count_208 + inc_207 - dec_207; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_207 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_207 <= count_207 + inc_206 - dec_206; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_206 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_206 <= count_206 + inc_205 - dec_205; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_205 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_205 <= count_205 + inc_204 - dec_204; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_204 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_204 <= count_204 + inc_203 - dec_203; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_203 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_203 <= count_203 + inc_202 - dec_202; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_202 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_202 <= count_202 + inc_201 - dec_201; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_201 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_201 <= count_201 + inc_200 - dec_200; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_200 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_200 <= count_200 + inc_199 - dec_199; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_199 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_199 <= count_199 + inc_198 - dec_198; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_198 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_198 <= count_198 + inc_197 - dec_197; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_197 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_197 <= count_197 + inc_196 - dec_196; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_196 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_196 <= count_196 + inc_195 - dec_195; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_195 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_195 <= count_195 + inc_194 - dec_194; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_194 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_194 <= count_194 + inc_193 - dec_193; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_193 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_193 <= count_193 + inc_192 - dec_192; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_192 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_192 <= count_192 + inc_191 - dec_191; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_191 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_191 <= count_191 + inc_190 - dec_190; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_190 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_190 <= count_190 + inc_189 - dec_189; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_189 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_189 <= count_189 + inc_188 - dec_188; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_188 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_188 <= count_188 + inc_187 - dec_187; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_187 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_187 <= count_187 + inc_186 - dec_186; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_186 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_186 <= count_186 + inc_185 - dec_185; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_185 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_185 <= count_185 + inc_184 - dec_184; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_184 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_184 <= count_184 + inc_183 - dec_183; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_183 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_183 <= count_183 + inc_182 - dec_182; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_182 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_182 <= count_182 + inc_181 - dec_181; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_181 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_181 <= count_181 + inc_180 - dec_180; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_180 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_180 <= count_180 + inc_179 - dec_179; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_179 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_179 <= count_179 + inc_178 - dec_178; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_178 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_178 <= count_178 + inc_177 - dec_177; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_177 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_177 <= count_177 + inc_176 - dec_176; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_176 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_176 <= count_176 + inc_175 - dec_175; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_175 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_175 <= count_175 + inc_174 - dec_174; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_174 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_174 <= count_174 + inc_173 - dec_173; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_173 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_173 <= count_173 + inc_172 - dec_172; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_172 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_172 <= count_172 + inc_171 - dec_171; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_171 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_171 <= count_171 + inc_170 - dec_170; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_170 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_170 <= count_170 + inc_169 - dec_169; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_169 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_169 <= count_169 + inc_168 - dec_168; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_168 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_168 <= count_168 + inc_167 - dec_167; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_167 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_167 <= count_167 + inc_166 - dec_166; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_166 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_166 <= count_166 + inc_165 - dec_165; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_165 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_165 <= count_165 + inc_164 - dec_164; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_164 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_164 <= count_164 + inc_163 - dec_163; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_163 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_163 <= count_163 + inc_162 - dec_162; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_162 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_162 <= count_162 + inc_161 - dec_161; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_161 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_161 <= count_161 + inc_160 - dec_160; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_160 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_160 <= count_160 + inc_159 - dec_159; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_159 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_159 <= count_159 + inc_158 - dec_158; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_158 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_158 <= count_158 + inc_157 - dec_157; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_157 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_157 <= count_157 + inc_156 - dec_156; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_156 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_156 <= count_156 + inc_155 - dec_155; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_155 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_155 <= count_155 + inc_154 - dec_154; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_154 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_154 <= count_154 + inc_153 - dec_153; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_153 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_153 <= count_153 + inc_152 - dec_152; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_152 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_152 <= count_152 + inc_151 - dec_151; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_151 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_151 <= count_151 + inc_150 - dec_150; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_150 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_150 <= count_150 + inc_149 - dec_149; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_149 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_149 <= count_149 + inc_148 - dec_148; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_148 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_148 <= count_148 + inc_147 - dec_147; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_147 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_147 <= count_147 + inc_146 - dec_146; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_146 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_146 <= count_146 + inc_145 - dec_145; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_145 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_145 <= count_145 + inc_144 - dec_144; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_144 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_144 <= count_144 + inc_143 - dec_143; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_143 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_143 <= count_143 + inc_142 - dec_142; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_142 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_142 <= count_142 + inc_141 - dec_141; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_141 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_141 <= count_141 + inc_140 - dec_140; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_140 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_140 <= count_140 + inc_139 - dec_139; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_139 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_139 <= count_139 + inc_138 - dec_138; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_138 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_138 <= count_138 + inc_137 - dec_137; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_137 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_137 <= count_137 + inc_136 - dec_136; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_136 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_136 <= count_136 + inc_135 - dec_135; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_135 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_135 <= count_135 + inc_134 - dec_134; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_134 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_134 <= count_134 + inc_133 - dec_133; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_133 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_133 <= count_133 + inc_132 - dec_132; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_132 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_132 <= count_132 + inc_131 - dec_131; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_131 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_131 <= count_131 + inc_130 - dec_130; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_130 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_130 <= count_130 + inc_129 - dec_129; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_129 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_129 <= count_129 + inc_128 - dec_128; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_128 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_128 <= count_128 + inc_127 - dec_127; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_127 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_127 <= count_127 + inc_126 - dec_126; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_126 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_126 <= count_126 + inc_125 - dec_125; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_125 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_125 <= count_125 + inc_124 - dec_124; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_124 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_124 <= count_124 + inc_123 - dec_123; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_123 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_123 <= count_123 + inc_122 - dec_122; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_122 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_122 <= count_122 + inc_121 - dec_121; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_121 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_121 <= count_121 + inc_120 - dec_120; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_120 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_120 <= count_120 + inc_119 - dec_119; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_119 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_119 <= count_119 + inc_118 - dec_118; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_118 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_118 <= count_118 + inc_117 - dec_117; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_117 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_117 <= count_117 + inc_116 - dec_116; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_116 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_116 <= count_116 + inc_115 - dec_115; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_115 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_115 <= count_115 + inc_114 - dec_114; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_114 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_114 <= count_114 + inc_113 - dec_113; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_113 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_113 <= count_113 + inc_112 - dec_112; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_112 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_112 <= count_112 + inc_111 - dec_111; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_111 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_111 <= count_111 + inc_110 - dec_110; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_110 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_110 <= count_110 + inc_109 - dec_109; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_109 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_109 <= count_109 + inc_108 - dec_108; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_108 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_108 <= count_108 + inc_107 - dec_107; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_107 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_107 <= count_107 + inc_106 - dec_106; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_106 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_106 <= count_106 + inc_105 - dec_105; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_105 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_105 <= count_105 + inc_104 - dec_104; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_104 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_104 <= count_104 + inc_103 - dec_103; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_103 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_103 <= count_103 + inc_102 - dec_102; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_102 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_102 <= count_102 + inc_101 - dec_101; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_101 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_101 <= count_101 + inc_100 - dec_100; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_100 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_100 <= count_100 + inc_99 - dec_99; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_99 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_99 <= count_99 + inc_98 - dec_98; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_98 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_98 <= count_98 + inc_97 - dec_97; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_97 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_97 <= count_97 + inc_96 - dec_96; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_96 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_96 <= count_96 + inc_95 - dec_95; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_95 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_95 <= count_95 + inc_94 - dec_94; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_94 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_94 <= count_94 + inc_93 - dec_93; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_93 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_93 <= count_93 + inc_92 - dec_92; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_92 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_92 <= count_92 + inc_91 - dec_91; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_91 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_91 <= count_91 + inc_90 - dec_90; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_90 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_90 <= count_90 + inc_89 - dec_89; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_89 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_89 <= count_89 + inc_88 - dec_88; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_88 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_88 <= count_88 + inc_87 - dec_87; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_87 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_87 <= count_87 + inc_86 - dec_86; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_86 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_86 <= count_86 + inc_85 - dec_85; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_85 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_85 <= count_85 + inc_84 - dec_84; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_84 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_84 <= count_84 + inc_83 - dec_83; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_83 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_83 <= count_83 + inc_82 - dec_82; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_82 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_82 <= count_82 + inc_81 - dec_81; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_81 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_81 <= count_81 + inc_80 - dec_80; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_80 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_80 <= count_80 + inc_79 - dec_79; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_79 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_79 <= count_79 + inc_78 - dec_78; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_78 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_78 <= count_78 + inc_77 - dec_77; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_77 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_77 <= count_77 + inc_76 - dec_76; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_76 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_76 <= count_76 + inc_75 - dec_75; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_75 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_75 <= count_75 + inc_74 - dec_74; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_74 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_74 <= count_74 + inc_73 - dec_73; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_73 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_73 <= count_73 + inc_72 - dec_72; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_72 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_72 <= count_72 + inc_71 - dec_71; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_71 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_71 <= count_71 + inc_70 - dec_70; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_70 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_70 <= count_70 + inc_69 - dec_69; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_69 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_69 <= count_69 + inc_68 - dec_68; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_68 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_68 <= count_68 + inc_67 - dec_67; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_67 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_67 <= count_67 + inc_66 - dec_66; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_66 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_66 <= count_66 + inc_65 - dec_65; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_65 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_65 <= count_65 + inc_64 - dec_64; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_64 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_64 <= count_64 + inc_63 - dec_63; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_63 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_63 <= count_63 + inc_62 - dec_62; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_62 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_62 <= count_62 + inc_61 - dec_61; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_61 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_61 <= count_61 + inc_60 - dec_60; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_60 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_60 <= count_60 + inc_59 - dec_59; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_59 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_59 <= count_59 + inc_58 - dec_58; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_58 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_58 <= count_58 + inc_57 - dec_57; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_57 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_57 <= count_57 + inc_56 - dec_56; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_56 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_56 <= count_56 + inc_55 - dec_55; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_55 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_55 <= count_55 + inc_54 - dec_54; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_54 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_54 <= count_54 + inc_53 - dec_53; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_53 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_53 <= count_53 + inc_52 - dec_52; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_52 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_52 <= count_52 + inc_51 - dec_51; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_51 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_51 <= count_51 + inc_50 - dec_50; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_50 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_50 <= count_50 + inc_49 - dec_49; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_49 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_49 <= count_49 + inc_48 - dec_48; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_48 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_48 <= count_48 + inc_47 - dec_47; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_47 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_47 <= count_47 + inc_46 - dec_46; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_46 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_46 <= count_46 + inc_45 - dec_45; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_45 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_45 <= count_45 + inc_44 - dec_44; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_44 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_44 <= count_44 + inc_43 - dec_43; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_43 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_43 <= count_43 + inc_42 - dec_42; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_42 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_42 <= count_42 + inc_41 - dec_41; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_41 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_41 <= count_41 + inc_40 - dec_40; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_40 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_40 <= count_40 + inc_39 - dec_39; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_39 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_39 <= count_39 + inc_38 - dec_38; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_38 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_38 <= count_38 + inc_37 - dec_37; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_37 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_37 <= count_37 + inc_36 - dec_36; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_36 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_36 <= count_36 + inc_35 - dec_35; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_35 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_35 <= count_35 + inc_34 - dec_34; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_34 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_34 <= count_34 + inc_33 - dec_33; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_33 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_33 <= count_33 + inc_32 - dec_32; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_32 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_32 <= count_32 + inc_31 - dec_31; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_31 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_31 <= count_31 + inc_30 - dec_30; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_30 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_30 <= count_30 + inc_29 - dec_29; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_29 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_29 <= count_29 + inc_28 - dec_28; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_28 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_28 <= count_28 + inc_27 - dec_27; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_27 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_27 <= count_27 + inc_26 - dec_26; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_26 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_26 <= count_26 + inc_25 - dec_25; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_25 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_25 <= count_25 + inc_24 - dec_24; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_24 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_24 <= count_24 + inc_23 - dec_23; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_23 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_23 <= count_23 + inc_22 - dec_22; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_22 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_22 <= count_22 + inc_21 - dec_21; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_21 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_21 <= count_21 + inc_20 - dec_20; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_20 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_20 <= count_20 + inc_19 - dec_19; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_19 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_19 <= count_19 + inc_18 - dec_18; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_18 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_18 <= count_18 + inc_17 - dec_17; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_17 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_17 <= count_17 + inc_16 - dec_16; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_16 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_16 <= count_16 + inc_15 - dec_15; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_15 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_15 <= count_15 + inc_14 - dec_14; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_14 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_14 <= count_14 + inc_13 - dec_13; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_13 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_13 <= count_13 + inc_12 - dec_12; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_12 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_12 <= count_12 + inc_11 - dec_11; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_11 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_11 <= count_11 + inc_10 - dec_10; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_10 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_10 <= count_10 + inc_9 - dec_9; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_9 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_9 <= count_9 + inc_8 - dec_8; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_8 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_8 <= count_8 + inc_7 - dec_7; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_7 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_7 <= count_7 + inc_6 - dec_6; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_6 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_6 <= count_6 + inc_5 - dec_5; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_5 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_5 <= count_5 + inc_4 - dec_4; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_4 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_4 <= count_4 + inc_3 - dec_3; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_3 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_3 <= count_3 + inc_2 - dec_2; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_2 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_2 <= count_2 + inc_1 - dec_1; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[ToAXI4.scala 254:28]
      count_1 <= 1'h0; // @[ToAXI4.scala 254:28]
    end else begin
      count_1 <= count_1 + inc - dec; // @[ToAXI4.scala 260:15]
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_T) begin
      if (a_first) begin
        if (a_isPut) begin
          counter <= beats1_decode;
        end else begin
          counter <= 3'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (reset) begin // @[ToAXI4.scala 161:30]
      doneAW <= 1'h0; // @[ToAXI4.scala 161:30]
    end else if (_T) begin
      doneAW <= ~a_last;
    end
    if (reset) begin // @[ToAXI4.scala 206:30]
      r_holds_d <= 1'h0; // @[ToAXI4.scala 206:30]
    end else if (_T_2) begin
      r_holds_d <= ~auto_out_r_bits_last;
    end
    if (auto_out_b_valid & ~bundleOut_0_b_ready) begin // @[ToAXI4.scala 210:42]
      b_delay <= _b_delay_T_1; // @[ToAXI4.scala 211:17]
    end else begin
      b_delay <= 3'h0; // @[ToAXI4.scala 213:17]
    end
    r_first <= reset | _GEN_1028; // @[ToAXI4.scala 224:{28,28}]
    if (r_first) begin // @[Reg.scala 17:18]
      r_denied_r <= _r_denied_T; // @[Reg.scala 17:22]
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec | count_1) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec | count_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc | idle) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc | idle)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_1 | count_2) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_1 | count_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_1 | idle_1) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_1 | idle_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_2 | count_3) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_2 | count_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_2 | idle_2) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_2 | idle_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_3 | count_4) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_3 | count_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_3 | idle_3) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_3 | idle_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_4 | count_5) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_4 | count_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_4 | idle_4) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_4 | idle_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_5 | count_6) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_5 | count_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_5 | idle_5) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_5 | idle_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_6 | count_7) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_6 | count_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_6 | idle_6) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_6 | idle_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_7 | count_8) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_7 | count_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_7 | idle_7) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_7 | idle_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_8 | count_9) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_8 | count_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_8 | idle_8) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_8 | idle_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_9 | count_10) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_9 | count_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_9 | idle_9) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_9 | idle_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_10 | count_11) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_10 | count_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_10 | idle_10) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_10 | idle_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_11 | count_12) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_11 | count_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_11 | idle_11) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_11 | idle_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_12 | count_13) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_12 | count_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_12 | idle_12) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_12 | idle_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_13 | count_14) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_13 | count_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_13 | idle_13) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_13 | idle_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_14 | count_15) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_14 | count_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_14 | idle_14) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_14 | idle_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_15 | count_16) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_15 | count_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_15 | idle_15) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_15 | idle_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_16 | count_17) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_16 | count_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_16 | idle_16) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_16 | idle_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_17 | count_18) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_17 | count_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_17 | idle_17) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_17 | idle_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_18 | count_19) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_18 | count_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_18 | idle_18) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_18 | idle_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_19 | count_20) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_19 | count_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_19 | idle_19) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_19 | idle_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_20 | count_21) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_20 | count_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_20 | idle_20) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_20 | idle_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_21 | count_22) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_21 | count_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_21 | idle_21) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_21 | idle_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_22 | count_23) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_22 | count_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_22 | idle_22) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_22 | idle_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_23 | count_24) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_23 | count_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_23 | idle_23) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_23 | idle_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_24 | count_25) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_24 | count_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_24 | idle_24) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_24 | idle_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_25 | count_26) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_25 | count_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_25 | idle_25) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_25 | idle_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_26 | count_27) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_26 | count_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_26 | idle_26) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_26 | idle_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_27 | count_28) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_27 | count_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_27 | idle_27) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_27 | idle_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_28 | count_29) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_28 | count_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_28 | idle_28) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_28 | idle_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_29 | count_30) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_29 | count_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_29 | idle_29) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_29 | idle_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_30 | count_31) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_30 | count_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_30 | idle_30) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_30 | idle_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_31 | count_32) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_31 | count_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_31 | idle_31) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_31 | idle_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_32 | count_33) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_32 | count_33)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_32 | idle_32) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_32 | idle_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_33 | count_34) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_33 | count_34)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_33 | idle_33) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_33 | idle_33)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_34 | count_35) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_34 | count_35)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_34 | idle_34) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_34 | idle_34)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_35 | count_36) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_35 | count_36)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_35 | idle_35) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_35 | idle_35)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_36 | count_37) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_36 | count_37)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_36 | idle_36) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_36 | idle_36)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_37 | count_38) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_37 | count_38)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_37 | idle_37) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_37 | idle_37)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_38 | count_39) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_38 | count_39)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_38 | idle_38) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_38 | idle_38)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_39 | count_40) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_39 | count_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_39 | idle_39) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_39 | idle_39)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_40 | count_41) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_40 | count_41)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_40 | idle_40) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_40 | idle_40)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_41 | count_42) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_41 | count_42)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_41 | idle_41) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_41 | idle_41)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_42 | count_43) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_42 | count_43)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_42 | idle_42) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_42 | idle_42)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_43 | count_44) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_43 | count_44)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_43 | idle_43) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_43 | idle_43)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_44 | count_45) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_44 | count_45)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_44 | idle_44) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_44 | idle_44)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_45 | count_46) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_45 | count_46)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_45 | idle_45) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_45 | idle_45)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_46 | count_47) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_46 | count_47)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_46 | idle_46) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_46 | idle_46)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_47 | count_48) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_47 | count_48)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_47 | idle_47) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_47 | idle_47)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_48 | count_49) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_48 | count_49)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_48 | idle_48) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_48 | idle_48)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_49 | count_50) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_49 | count_50)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_49 | idle_49) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_49 | idle_49)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_50 | count_51) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_50 | count_51)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_50 | idle_50) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_50 | idle_50)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_51 | count_52) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_51 | count_52)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_51 | idle_51) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_51 | idle_51)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_52 | count_53) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_52 | count_53)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_52 | idle_52) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_52 | idle_52)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_53 | count_54) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_53 | count_54)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_53 | idle_53) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_53 | idle_53)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_54 | count_55) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_54 | count_55)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_54 | idle_54) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_54 | idle_54)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_55 | count_56) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_55 | count_56)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_55 | idle_55) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_55 | idle_55)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_56 | count_57) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_56 | count_57)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_56 | idle_56) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_56 | idle_56)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_57 | count_58) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_57 | count_58)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_57 | idle_57) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_57 | idle_57)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_58 | count_59) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_58 | count_59)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_58 | idle_58) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_58 | idle_58)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_59 | count_60) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_59 | count_60)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_59 | idle_59) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_59 | idle_59)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_60 | count_61) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_60 | count_61)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_60 | idle_60) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_60 | idle_60)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_61 | count_62) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_61 | count_62)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_61 | idle_61) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_61 | idle_61)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_62 | count_63) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_62 | count_63)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_62 | idle_62) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_62 | idle_62)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_63 | count_64) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_63 | count_64)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_63 | idle_63) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_63 | idle_63)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_64 | count_65) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_64 | count_65)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_64 | idle_64) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_64 | idle_64)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_65 | count_66) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_65 | count_66)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_65 | idle_65) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_65 | idle_65)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_66 | count_67) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_66 | count_67)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_66 | idle_66) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_66 | idle_66)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_67 | count_68) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_67 | count_68)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_67 | idle_67) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_67 | idle_67)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_68 | count_69) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_68 | count_69)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_68 | idle_68) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_68 | idle_68)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_69 | count_70) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_69 | count_70)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_69 | idle_69) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_69 | idle_69)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_70 | count_71) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_70 | count_71)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_70 | idle_70) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_70 | idle_70)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_71 | count_72) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_71 | count_72)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_71 | idle_71) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_71 | idle_71)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_72 | count_73) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_72 | count_73)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_72 | idle_72) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_72 | idle_72)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_73 | count_74) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_73 | count_74)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_73 | idle_73) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_73 | idle_73)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_74 | count_75) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_74 | count_75)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_74 | idle_74) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_74 | idle_74)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_75 | count_76) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_75 | count_76)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_75 | idle_75) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_75 | idle_75)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_76 | count_77) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_76 | count_77)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_76 | idle_76) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_76 | idle_76)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_77 | count_78) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_77 | count_78)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_77 | idle_77) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_77 | idle_77)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_78 | count_79) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_78 | count_79)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_78 | idle_78) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_78 | idle_78)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_79 | count_80) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_79 | count_80)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_79 | idle_79) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_79 | idle_79)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_80 | count_81) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_80 | count_81)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_80 | idle_80) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_80 | idle_80)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_81 | count_82) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_81 | count_82)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_81 | idle_81) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_81 | idle_81)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_82 | count_83) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_82 | count_83)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_82 | idle_82) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_82 | idle_82)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_83 | count_84) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_83 | count_84)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_83 | idle_83) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_83 | idle_83)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_84 | count_85) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_84 | count_85)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_84 | idle_84) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_84 | idle_84)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_85 | count_86) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_85 | count_86)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_85 | idle_85) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_85 | idle_85)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_86 | count_87) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_86 | count_87)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_86 | idle_86) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_86 | idle_86)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_87 | count_88) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_87 | count_88)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_87 | idle_87) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_87 | idle_87)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_88 | count_89) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_88 | count_89)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_88 | idle_88) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_88 | idle_88)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_89 | count_90) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_89 | count_90)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_89 | idle_89) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_89 | idle_89)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_90 | count_91) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_90 | count_91)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_90 | idle_90) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_90 | idle_90)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_91 | count_92) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_91 | count_92)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_91 | idle_91) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_91 | idle_91)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_92 | count_93) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_92 | count_93)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_92 | idle_92) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_92 | idle_92)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_93 | count_94) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_93 | count_94)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_93 | idle_93) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_93 | idle_93)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_94 | count_95) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_94 | count_95)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_94 | idle_94) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_94 | idle_94)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_95 | count_96) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_95 | count_96)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_95 | idle_95) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_95 | idle_95)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_96 | count_97) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_96 | count_97)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_96 | idle_96) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_96 | idle_96)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_97 | count_98) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_97 | count_98)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_97 | idle_97) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_97 | idle_97)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_98 | count_99) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_98 | count_99)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_98 | idle_98) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_98 | idle_98)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_99 | count_100) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_99 | count_100)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_99 | idle_99) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_99 | idle_99)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_100 | count_101) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_100 | count_101)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_100 | idle_100) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_100 | idle_100)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_101 | count_102) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_101 | count_102)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_101 | idle_101) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_101 | idle_101)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_102 | count_103) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_102 | count_103)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_102 | idle_102) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_102 | idle_102)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_103 | count_104) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_103 | count_104)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_103 | idle_103) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_103 | idle_103)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_104 | count_105) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_104 | count_105)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_104 | idle_104) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_104 | idle_104)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_105 | count_106) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_105 | count_106)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_105 | idle_105) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_105 | idle_105)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_106 | count_107) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_106 | count_107)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_106 | idle_106) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_106 | idle_106)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_107 | count_108) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_107 | count_108)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_107 | idle_107) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_107 | idle_107)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_108 | count_109) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_108 | count_109)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_108 | idle_108) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_108 | idle_108)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_109 | count_110) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_109 | count_110)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_109 | idle_109) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_109 | idle_109)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_110 | count_111) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_110 | count_111)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_110 | idle_110) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_110 | idle_110)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_111 | count_112) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_111 | count_112)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_111 | idle_111) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_111 | idle_111)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_112 | count_113) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_112 | count_113)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_112 | idle_112) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_112 | idle_112)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_113 | count_114) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_113 | count_114)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_113 | idle_113) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_113 | idle_113)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_114 | count_115) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_114 | count_115)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_114 | idle_114) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_114 | idle_114)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_115 | count_116) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_115 | count_116)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_115 | idle_115) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_115 | idle_115)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_116 | count_117) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_116 | count_117)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_116 | idle_116) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_116 | idle_116)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_117 | count_118) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_117 | count_118)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_117 | idle_117) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_117 | idle_117)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_118 | count_119) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_118 | count_119)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_118 | idle_118) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_118 | idle_118)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_119 | count_120) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_119 | count_120)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_119 | idle_119) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_119 | idle_119)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_120 | count_121) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_120 | count_121)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_120 | idle_120) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_120 | idle_120)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_121 | count_122) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_121 | count_122)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_121 | idle_121) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_121 | idle_121)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_122 | count_123) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_122 | count_123)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_122 | idle_122) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_122 | idle_122)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_123 | count_124) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_123 | count_124)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_123 | idle_123) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_123 | idle_123)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_124 | count_125) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_124 | count_125)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_124 | idle_124) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_124 | idle_124)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_125 | count_126) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_125 | count_126)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_125 | idle_125) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_125 | idle_125)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_126 | count_127) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_126 | count_127)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_126 | idle_126) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_126 | idle_126)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_127 | count_128) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_127 | count_128)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_127 | idle_127) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_127 | idle_127)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_128 | count_129) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_128 | count_129)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_128 | idle_128) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_128 | idle_128)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_129 | count_130) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_129 | count_130)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_129 | idle_129) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_129 | idle_129)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_130 | count_131) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_130 | count_131)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_130 | idle_130) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_130 | idle_130)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_131 | count_132) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_131 | count_132)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_131 | idle_131) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_131 | idle_131)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_132 | count_133) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_132 | count_133)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_132 | idle_132) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_132 | idle_132)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_133 | count_134) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_133 | count_134)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_133 | idle_133) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_133 | idle_133)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_134 | count_135) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_134 | count_135)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_134 | idle_134) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_134 | idle_134)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_135 | count_136) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_135 | count_136)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_135 | idle_135) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_135 | idle_135)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_136 | count_137) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_136 | count_137)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_136 | idle_136) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_136 | idle_136)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_137 | count_138) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_137 | count_138)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_137 | idle_137) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_137 | idle_137)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_138 | count_139) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_138 | count_139)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_138 | idle_138) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_138 | idle_138)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_139 | count_140) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_139 | count_140)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_139 | idle_139) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_139 | idle_139)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_140 | count_141) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_140 | count_141)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_140 | idle_140) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_140 | idle_140)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_141 | count_142) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_141 | count_142)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_141 | idle_141) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_141 | idle_141)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_142 | count_143) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_142 | count_143)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_142 | idle_142) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_142 | idle_142)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_143 | count_144) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_143 | count_144)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_143 | idle_143) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_143 | idle_143)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_144 | count_145) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_144 | count_145)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_144 | idle_144) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_144 | idle_144)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_145 | count_146) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_145 | count_146)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_145 | idle_145) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_145 | idle_145)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_146 | count_147) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_146 | count_147)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_146 | idle_146) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_146 | idle_146)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_147 | count_148) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_147 | count_148)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_147 | idle_147) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_147 | idle_147)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_148 | count_149) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_148 | count_149)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_148 | idle_148) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_148 | idle_148)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_149 | count_150) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_149 | count_150)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_149 | idle_149) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_149 | idle_149)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_150 | count_151) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_150 | count_151)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_150 | idle_150) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_150 | idle_150)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_151 | count_152) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_151 | count_152)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_151 | idle_151) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_151 | idle_151)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_152 | count_153) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_152 | count_153)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_152 | idle_152) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_152 | idle_152)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_153 | count_154) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_153 | count_154)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_153 | idle_153) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_153 | idle_153)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_154 | count_155) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_154 | count_155)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_154 | idle_154) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_154 | idle_154)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_155 | count_156) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_155 | count_156)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_155 | idle_155) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_155 | idle_155)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_156 | count_157) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_156 | count_157)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_156 | idle_156) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_156 | idle_156)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_157 | count_158) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_157 | count_158)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_157 | idle_157) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_157 | idle_157)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_158 | count_159) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_158 | count_159)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_158 | idle_158) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_158 | idle_158)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_159 | count_160) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_159 | count_160)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_159 | idle_159) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_159 | idle_159)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_160 | count_161) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_160 | count_161)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_160 | idle_160) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_160 | idle_160)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_161 | count_162) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_161 | count_162)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_161 | idle_161) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_161 | idle_161)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_162 | count_163) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_162 | count_163)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_162 | idle_162) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_162 | idle_162)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_163 | count_164) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_163 | count_164)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_163 | idle_163) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_163 | idle_163)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_164 | count_165) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_164 | count_165)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_164 | idle_164) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_164 | idle_164)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_165 | count_166) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_165 | count_166)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_165 | idle_165) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_165 | idle_165)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_166 | count_167) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_166 | count_167)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_166 | idle_166) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_166 | idle_166)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_167 | count_168) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_167 | count_168)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_167 | idle_167) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_167 | idle_167)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_168 | count_169) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_168 | count_169)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_168 | idle_168) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_168 | idle_168)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_169 | count_170) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_169 | count_170)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_169 | idle_169) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_169 | idle_169)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_170 | count_171) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_170 | count_171)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_170 | idle_170) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_170 | idle_170)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_171 | count_172) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_171 | count_172)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_171 | idle_171) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_171 | idle_171)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_172 | count_173) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_172 | count_173)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_172 | idle_172) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_172 | idle_172)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_173 | count_174) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_173 | count_174)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_173 | idle_173) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_173 | idle_173)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_174 | count_175) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_174 | count_175)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_174 | idle_174) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_174 | idle_174)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_175 | count_176) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_175 | count_176)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_175 | idle_175) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_175 | idle_175)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_176 | count_177) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_176 | count_177)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_176 | idle_176) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_176 | idle_176)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_177 | count_178) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_177 | count_178)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_177 | idle_177) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_177 | idle_177)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_178 | count_179) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_178 | count_179)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_178 | idle_178) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_178 | idle_178)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_179 | count_180) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_179 | count_180)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_179 | idle_179) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_179 | idle_179)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_180 | count_181) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_180 | count_181)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_180 | idle_180) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_180 | idle_180)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_181 | count_182) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_181 | count_182)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_181 | idle_181) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_181 | idle_181)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_182 | count_183) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_182 | count_183)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_182 | idle_182) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_182 | idle_182)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_183 | count_184) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_183 | count_184)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_183 | idle_183) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_183 | idle_183)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_184 | count_185) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_184 | count_185)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_184 | idle_184) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_184 | idle_184)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_185 | count_186) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_185 | count_186)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_185 | idle_185) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_185 | idle_185)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_186 | count_187) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_186 | count_187)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_186 | idle_186) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_186 | idle_186)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_187 | count_188) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_187 | count_188)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_187 | idle_187) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_187 | idle_187)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_188 | count_189) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_188 | count_189)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_188 | idle_188) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_188 | idle_188)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_189 | count_190) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_189 | count_190)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_189 | idle_189) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_189 | idle_189)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_190 | count_191) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_190 | count_191)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_190 | idle_190) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_190 | idle_190)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_191 | count_192) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_191 | count_192)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_191 | idle_191) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_191 | idle_191)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_192 | count_193) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_192 | count_193)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_192 | idle_192) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_192 | idle_192)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_193 | count_194) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_193 | count_194)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_193 | idle_193) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_193 | idle_193)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_194 | count_195) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_194 | count_195)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_194 | idle_194) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_194 | idle_194)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_195 | count_196) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_195 | count_196)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_195 | idle_195) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_195 | idle_195)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_196 | count_197) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_196 | count_197)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_196 | idle_196) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_196 | idle_196)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_197 | count_198) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_197 | count_198)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_197 | idle_197) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_197 | idle_197)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_198 | count_199) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_198 | count_199)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_198 | idle_198) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_198 | idle_198)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_199 | count_200) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_199 | count_200)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_199 | idle_199) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_199 | idle_199)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_200 | count_201) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_200 | count_201)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_200 | idle_200) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_200 | idle_200)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_201 | count_202) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_201 | count_202)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_201 | idle_201) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_201 | idle_201)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_202 | count_203) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_202 | count_203)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_202 | idle_202) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_202 | idle_202)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_203 | count_204) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_203 | count_204)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_203 | idle_203) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_203 | idle_203)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_204 | count_205) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_204 | count_205)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_204 | idle_204) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_204 | idle_204)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_205 | count_206) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_205 | count_206)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_205 | idle_205) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_205 | idle_205)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_206 | count_207) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_206 | count_207)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_206 | idle_206) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_206 | idle_206)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_207 | count_208) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_207 | count_208)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_207 | idle_207) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_207 | idle_207)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_208 | count_209) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_208 | count_209)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_208 | idle_208) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_208 | idle_208)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_209 | count_210) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_209 | count_210)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_209 | idle_209) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_209 | idle_209)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_210 | count_211) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_210 | count_211)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_210 | idle_210) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_210 | idle_210)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_211 | count_212) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_211 | count_212)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_211 | idle_211) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_211 | idle_211)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_212 | count_213) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_212 | count_213)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_212 | idle_212) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_212 | idle_212)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_213 | count_214) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_213 | count_214)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_213 | idle_213) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_213 | idle_213)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_214 | count_215) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_214 | count_215)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_214 | idle_214) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_214 | idle_214)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_215 | count_216) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_215 | count_216)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_215 | idle_215) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_215 | idle_215)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_216 | count_217) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_216 | count_217)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_216 | idle_216) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_216 | idle_216)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_217 | count_218) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_217 | count_218)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_217 | idle_217) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_217 | idle_217)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_218 | count_219) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_218 | count_219)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_218 | idle_218) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_218 | idle_218)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_219 | count_220) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_219 | count_220)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_219 | idle_219) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_219 | idle_219)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_220 | count_221) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_220 | count_221)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_220 | idle_220) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_220 | idle_220)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_221 | count_222) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_221 | count_222)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_221 | idle_221) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_221 | idle_221)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_222 | count_223) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_222 | count_223)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_222 | idle_222) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_222 | idle_222)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_223 | count_224) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_223 | count_224)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_223 | idle_223) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_223 | idle_223)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_224 | count_225) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_224 | count_225)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_224 | idle_224) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_224 | idle_224)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_225 | count_226) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_225 | count_226)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_225 | idle_225) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_225 | idle_225)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_226 | count_227) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_226 | count_227)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_226 | idle_226) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_226 | idle_226)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_227 | count_228) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_227 | count_228)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_227 | idle_227) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_227 | idle_227)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_228 | count_229) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_228 | count_229)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_228 | idle_228) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_228 | idle_228)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_229 | count_230) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_229 | count_230)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_229 | idle_229) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_229 | idle_229)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_230 | count_231) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_230 | count_231)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_230 | idle_230) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_230 | idle_230)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_231 | count_232) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_231 | count_232)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_231 | idle_231) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_231 | idle_231)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_232 | count_233) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_232 | count_233)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_232 | idle_232) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_232 | idle_232)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_233 | count_234) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_233 | count_234)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_233 | idle_233) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_233 | idle_233)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_234 | count_235) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_234 | count_235)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_234 | idle_234) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_234 | idle_234)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_235 | count_236) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_235 | count_236)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_235 | idle_235) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_235 | idle_235)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_236 | count_237) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_236 | count_237)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_236 | idle_236) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_236 | idle_236)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_237 | count_238) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_237 | count_238)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_237 | idle_237) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_237 | idle_237)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_238 | count_239) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_238 | count_239)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_238 | idle_238) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_238 | idle_238)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_239 | count_240) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_239 | count_240)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_239 | idle_239) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_239 | idle_239)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_240 | count_241) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_240 | count_241)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_240 | idle_240) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_240 | idle_240)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_241 | count_242) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_241 | count_242)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_241 | idle_241) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_241 | idle_241)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_242 | count_243) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_242 | count_243)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_242 | idle_242) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_242 | idle_242)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_243 | count_244) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_243 | count_244)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_243 | idle_243) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_243 | idle_243)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_244 | count_245) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_244 | count_245)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_244 | idle_244) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_244 | idle_244)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_245 | count_246) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_245 | count_246)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_245 | idle_245) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_245 | idle_245)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_246 | count_247) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_246 | count_247)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_246 | idle_246) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_246 | idle_246)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_247 | count_248) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_247 | count_248)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_247 | idle_247) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_247 | idle_247)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_248 | count_249) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_248 | count_249)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_248 | idle_248) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_248 | idle_248)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_249 | count_250) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_249 | count_250)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_249 | idle_249) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_249 | idle_249)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_250 | count_251) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_250 | count_251)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_250 | idle_250) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_250 | idle_250)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_251 | count_252) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_251 | count_252)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_251 | idle_251) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_251 | idle_251)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_252 | count_253) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_252 | count_253)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_252 | idle_252) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_252 | idle_252)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_253 | count_254) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_253 | count_254)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_253 | idle_253) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_253 | idle_253)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_254 | count_255) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_254 | count_255)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_254 | idle_254) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_254 | idle_254)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_255 | count_256) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_255 | count_256)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_255 | idle_255) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_255 | idle_255)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_256 | count_257) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_256 | count_257)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_256 | idle_256) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_256 | idle_256)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_257 | count_258) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_257 | count_258)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_257 | idle_257) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_257 | idle_257)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_258 | count_259) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_258 | count_259)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_258 | idle_258) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_258 | idle_258)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_259 | count_260) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_259 | count_260)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_259 | idle_259) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_259 | idle_259)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_260 | count_261) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_260 | count_261)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_260 | idle_260) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_260 | idle_260)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_261 | count_262) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_261 | count_262)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_261 | idle_261) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_261 | idle_261)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_262 | count_263) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_262 | count_263)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_262 | idle_262) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_262 | idle_262)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_263 | count_264) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_263 | count_264)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_263 | idle_263) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_263 | idle_263)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_264 | count_265) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_264 | count_265)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_264 | idle_264) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_264 | idle_264)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_265 | count_266) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_265 | count_266)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_265 | idle_265) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_265 | idle_265)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_266 | count_267) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_266 | count_267)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_266 | idle_266) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_266 | idle_266)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_267 | count_268) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_267 | count_268)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_267 | idle_267) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_267 | idle_267)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_268 | count_269) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_268 | count_269)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_268 | idle_268) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_268 | idle_268)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_269 | count_270) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_269 | count_270)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_269 | idle_269) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_269 | idle_269)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_270 | count_271) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_270 | count_271)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_270 | idle_270) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_270 | idle_270)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_271 | count_272) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_271 | count_272)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_271 | idle_271) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_271 | idle_271)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_272 | count_273) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_272 | count_273)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_272 | idle_272) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_272 | idle_272)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_273 | count_274) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_273 | count_274)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_273 | idle_273) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_273 | idle_273)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_274 | count_275) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_274 | count_275)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_274 | idle_274) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_274 | idle_274)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_275 | count_276) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_275 | count_276)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_275 | idle_275) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_275 | idle_275)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_276 | count_277) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_276 | count_277)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_276 | idle_276) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_276 | idle_276)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_277 | count_278) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_277 | count_278)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_277 | idle_277) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_277 | idle_277)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_278 | count_279) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_278 | count_279)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_278 | idle_278) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_278 | idle_278)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_279 | count_280) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_279 | count_280)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_279 | idle_279) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_279 | idle_279)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_280 | count_281) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_280 | count_281)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_280 | idle_280) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_280 | idle_280)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_281 | count_282) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_281 | count_282)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_281 | idle_281) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_281 | idle_281)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_282 | count_283) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_282 | count_283)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_282 | idle_282) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_282 | idle_282)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_283 | count_284) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_283 | count_284)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_283 | idle_283) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_283 | idle_283)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_284 | count_285) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_284 | count_285)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_284 | idle_284) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_284 | idle_284)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_285 | count_286) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_285 | count_286)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_285 | idle_285) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_285 | idle_285)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_286 | count_287) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_286 | count_287)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_286 | idle_286) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_286 | idle_286)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_287 | count_288) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_287 | count_288)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_287 | idle_287) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_287 | idle_287)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_288 | count_289) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_288 | count_289)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_288 | idle_288) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_288 | idle_288)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_289 | count_290) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_289 | count_290)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_289 | idle_289) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_289 | idle_289)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_290 | count_291) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_290 | count_291)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_290 | idle_290) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_290 | idle_290)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_291 | count_292) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_291 | count_292)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_291 | idle_291) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_291 | idle_291)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_292 | count_293) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_292 | count_293)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_292 | idle_292) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_292 | idle_292)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_293 | count_294) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_293 | count_294)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_293 | idle_293) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_293 | idle_293)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_294 | count_295) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_294 | count_295)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_294 | idle_294) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_294 | idle_294)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_295 | count_296) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_295 | count_296)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_295 | idle_295) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_295 | idle_295)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_296 | count_297) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_296 | count_297)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_296 | idle_296) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_296 | idle_296)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_297 | count_298) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_297 | count_298)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_297 | idle_297) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_297 | idle_297)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_298 | count_299) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_298 | count_299)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_298 | idle_298) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_298 | idle_298)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_299 | count_300) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_299 | count_300)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_299 | idle_299) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_299 | idle_299)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_300 | count_301) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_300 | count_301)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_300 | idle_300) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_300 | idle_300)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_301 | count_302) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_301 | count_302)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_301 | idle_301) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_301 | idle_301)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_302 | count_303) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_302 | count_303)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_302 | idle_302) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_302 | idle_302)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_303 | count_304) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_303 | count_304)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_303 | idle_303) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_303 | idle_303)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_304 | count_305) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_304 | count_305)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_304 | idle_304) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_304 | idle_304)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_305 | count_306) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_305 | count_306)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_305 | idle_305) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_305 | idle_305)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_306 | count_307) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_306 | count_307)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_306 | idle_306) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_306 | idle_306)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_307 | count_308) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_307 | count_308)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_307 | idle_307) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_307 | idle_307)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_308 | count_309) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_308 | count_309)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_308 | idle_308) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_308 | idle_308)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_309 | count_310) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_309 | count_310)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_309 | idle_309) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_309 | idle_309)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_310 | count_311) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_310 | count_311)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_310 | idle_310) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_310 | idle_310)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_311 | count_312) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_311 | count_312)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_311 | idle_311) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_311 | idle_311)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_312 | count_313) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_312 | count_313)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_312 | idle_312) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_312 | idle_312)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_313 | count_314) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_313 | count_314)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_313 | idle_313) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_313 | idle_313)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_314 | count_315) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_314 | count_315)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_314 | idle_314) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_314 | idle_314)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_315 | count_316) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_315 | count_316)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_315 | idle_315) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_315 | idle_315)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_316 | count_317) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_316 | count_317)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_316 | idle_316) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_316 | idle_316)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_317 | count_318) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_317 | count_318)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_317 | idle_317) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_317 | idle_317)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_318 | count_319) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_318 | count_319)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_318 | idle_318) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_318 | idle_318)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_319 | count_320) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_319 | count_320)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_319 | idle_319) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_319 | idle_319)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_320 | count_321) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_320 | count_321)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_320 | idle_320) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_320 | idle_320)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_321 | count_322) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_321 | count_322)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_321 | idle_321) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_321 | idle_321)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_322 | count_323) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_322 | count_323)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_322 | idle_322) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_322 | idle_322)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_323 | count_324) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_323 | count_324)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_323 | idle_323) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_323 | idle_323)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_324 | count_325) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_324 | count_325)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_324 | idle_324) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_324 | idle_324)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_325 | count_326) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_325 | count_326)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_325 | idle_325) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_325 | idle_325)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_326 | count_327) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_326 | count_327)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_326 | idle_326) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_326 | idle_326)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_327 | count_328) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_327 | count_328)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_327 | idle_327) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_327 | idle_327)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_328 | count_329) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_328 | count_329)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_328 | idle_328) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_328 | idle_328)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_329 | count_330) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_329 | count_330)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_329 | idle_329) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_329 | idle_329)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_330 | count_331) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_330 | count_331)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_330 | idle_330) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_330 | idle_330)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_331 | count_332) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_331 | count_332)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_331 | idle_331) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_331 | idle_331)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_332 | count_333) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_332 | count_333)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_332 | idle_332) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_332 | idle_332)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_333 | count_334) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_333 | count_334)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_333 | idle_333) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_333 | idle_333)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_334 | count_335) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_334 | count_335)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_334 | idle_334) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_334 | idle_334)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_335 | count_336) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_335 | count_336)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_335 | idle_335) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_335 | idle_335)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_336 | count_337) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_336 | count_337)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_336 | idle_336) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_336 | idle_336)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_337 | count_338) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_337 | count_338)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_337 | idle_337) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_337 | idle_337)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_338 | count_339) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_338 | count_339)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_338 | idle_338) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_338 | idle_338)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_339 | count_340) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_339 | count_340)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_339 | idle_339) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_339 | idle_339)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_340 | count_341) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_340 | count_341)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_340 | idle_340) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_340 | idle_340)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_341 | count_342) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_341 | count_342)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_341 | idle_341) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_341 | idle_341)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_342 | count_343) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_342 | count_343)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_342 | idle_342) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_342 | idle_342)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_343 | count_344) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_343 | count_344)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_343 | idle_343) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_343 | idle_343)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_344 | count_345) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_344 | count_345)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_344 | idle_344) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_344 | idle_344)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_345 | count_346) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_345 | count_346)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_345 | idle_345) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_345 | idle_345)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_346 | count_347) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_346 | count_347)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_346 | idle_346) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_346 | idle_346)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_347 | count_348) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_347 | count_348)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_347 | idle_347) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_347 | idle_347)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_348 | count_349) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_348 | count_349)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_348 | idle_348) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_348 | idle_348)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_349 | count_350) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_349 | count_350)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_349 | idle_349) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_349 | idle_349)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_350 | count_351) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_350 | count_351)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_350 | idle_350) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_350 | idle_350)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_351 | count_352) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_351 | count_352)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_351 | idle_351) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_351 | idle_351)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_352 | count_353) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_352 | count_353)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_352 | idle_352) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_352 | idle_352)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_353 | count_354) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_353 | count_354)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_353 | idle_353) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_353 | idle_353)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_354 | count_355) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_354 | count_355)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_354 | idle_354) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_354 | idle_354)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_355 | count_356) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_355 | count_356)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_355 | idle_355) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_355 | idle_355)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_356 | count_357) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_356 | count_357)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_356 | idle_356) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_356 | idle_356)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_357 | count_358) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_357 | count_358)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_357 | idle_357) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_357 | idle_357)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_358 | count_359) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_358 | count_359)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_358 | idle_358) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_358 | idle_358)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_359 | count_360) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_359 | count_360)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_359 | idle_359) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_359 | idle_359)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_360 | count_361) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_360 | count_361)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_360 | idle_360) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_360 | idle_360)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_361 | count_362) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_361 | count_362)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_361 | idle_361) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_361 | idle_361)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_362 | count_363) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_362 | count_363)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_362 | idle_362) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_362 | idle_362)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_363 | count_364) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_363 | count_364)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_363 | idle_363) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_363 | idle_363)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_364 | count_365) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_364 | count_365)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_364 | idle_364) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_364 | idle_364)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_365 | count_366) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_365 | count_366)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_365 | idle_365) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_365 | idle_365)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_366 | count_367) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_366 | count_367)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_366 | idle_366) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_366 | idle_366)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_367 | count_368) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_367 | count_368)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_367 | idle_367) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_367 | idle_367)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_368 | count_369) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_368 | count_369)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_368 | idle_368) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_368 | idle_368)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_369 | count_370) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_369 | count_370)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_369 | idle_369) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_369 | idle_369)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_370 | count_371) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_370 | count_371)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_370 | idle_370) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_370 | idle_370)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_371 | count_372) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_371 | count_372)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_371 | idle_371) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_371 | idle_371)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_372 | count_373) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_372 | count_373)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_372 | idle_372) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_372 | idle_372)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_373 | count_374) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_373 | count_374)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_373 | idle_373) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_373 | idle_373)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_374 | count_375) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_374 | count_375)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_374 | idle_374) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_374 | idle_374)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_375 | count_376) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_375 | count_376)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_375 | idle_375) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_375 | idle_375)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_376 | count_377) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_376 | count_377)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_376 | idle_376) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_376 | idle_376)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_377 | count_378) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_377 | count_378)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_377 | idle_377) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_377 | idle_377)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_378 | count_379) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_378 | count_379)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_378 | idle_378) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_378 | idle_378)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_379 | count_380) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_379 | count_380)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_379 | idle_379) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_379 | idle_379)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_380 | count_381) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_380 | count_381)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_380 | idle_380) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_380 | idle_380)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_381 | count_382) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_381 | count_382)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_381 | idle_381) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_381 | idle_381)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_382 | count_383) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_382 | count_383)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_382 | idle_382) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_382 | idle_382)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_383 | count_384) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_383 | count_384)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_383 | idle_383) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_383 | idle_383)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_384 | count_385) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_384 | count_385)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_384 | idle_384) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_384 | idle_384)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_385 | count_386) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_385 | count_386)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_385 | idle_385) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_385 | idle_385)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_386 | count_387) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_386 | count_387)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_386 | idle_386) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_386 | idle_386)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_387 | count_388) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_387 | count_388)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_387 | idle_387) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_387 | idle_387)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_388 | count_389) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_388 | count_389)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_388 | idle_388) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_388 | idle_388)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_389 | count_390) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_389 | count_390)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_389 | idle_389) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_389 | idle_389)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_390 | count_391) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_390 | count_391)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_390 | idle_390) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_390 | idle_390)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_391 | count_392) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_391 | count_392)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_391 | idle_391) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_391 | idle_391)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_392 | count_393) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_392 | count_393)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_392 | idle_392) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_392 | idle_392)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_393 | count_394) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_393 | count_394)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_393 | idle_393) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_393 | idle_393)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_394 | count_395) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_394 | count_395)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_394 | idle_394) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_394 | idle_394)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_395 | count_396) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_395 | count_396)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_395 | idle_395) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_395 | idle_395)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_396 | count_397) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_396 | count_397)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_396 | idle_396) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_396 | idle_396)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_397 | count_398) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_397 | count_398)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_397 | idle_397) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_397 | idle_397)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_398 | count_399) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_398 | count_399)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_398 | idle_398) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_398 | idle_398)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_399 | count_400) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_399 | count_400)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_399 | idle_399) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_399 | idle_399)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_400 | count_401) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_400 | count_401)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_400 | idle_400) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_400 | idle_400)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_401 | count_402) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_401 | count_402)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_401 | idle_401) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_401 | idle_401)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_402 | count_403) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_402 | count_403)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_402 | idle_402) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_402 | idle_402)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_403 | count_404) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_403 | count_404)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_403 | idle_403) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_403 | idle_403)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_404 | count_405) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_404 | count_405)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_404 | idle_404) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_404 | idle_404)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_405 | count_406) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_405 | count_406)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_405 | idle_405) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_405 | idle_405)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_406 | count_407) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_406 | count_407)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_406 | idle_406) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_406 | idle_406)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_407 | count_408) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_407 | count_408)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_407 | idle_407) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_407 | idle_407)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_408 | count_409) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_408 | count_409)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_408 | idle_408) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_408 | idle_408)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_409 | count_410) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_409 | count_410)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_409 | idle_409) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_409 | idle_409)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_410 | count_411) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_410 | count_411)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_410 | idle_410) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_410 | idle_410)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_411 | count_412) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_411 | count_412)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_411 | idle_411) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_411 | idle_411)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_412 | count_413) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_412 | count_413)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_412 | idle_412) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_412 | idle_412)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_413 | count_414) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_413 | count_414)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_413 | idle_413) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_413 | idle_413)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_414 | count_415) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_414 | count_415)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_414 | idle_414) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_414 | idle_414)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_415 | count_416) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_415 | count_416)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_415 | idle_415) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_415 | idle_415)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_416 | count_417) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_416 | count_417)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_416 | idle_416) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_416 | idle_416)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_417 | count_418) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_417 | count_418)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_417 | idle_417) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_417 | idle_417)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_418 | count_419) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_418 | count_419)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_418 | idle_418) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_418 | idle_418)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_419 | count_420) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_419 | count_420)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_419 | idle_419) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_419 | idle_419)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_420 | count_421) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_420 | count_421)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_420 | idle_420) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_420 | idle_420)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_421 | count_422) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_421 | count_422)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_421 | idle_421) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_421 | idle_421)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_422 | count_423) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_422 | count_423)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_422 | idle_422) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_422 | idle_422)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_423 | count_424) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_423 | count_424)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_423 | idle_423) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_423 | idle_423)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_424 | count_425) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_424 | count_425)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_424 | idle_424) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_424 | idle_424)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_425 | count_426) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_425 | count_426)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_425 | idle_425) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_425 | idle_425)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_426 | count_427) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_426 | count_427)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_426 | idle_426) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_426 | idle_426)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_427 | count_428) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_427 | count_428)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_427 | idle_427) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_427 | idle_427)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_428 | count_429) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_428 | count_429)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_428 | idle_428) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_428 | idle_428)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_429 | count_430) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_429 | count_430)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_429 | idle_429) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_429 | idle_429)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_430 | count_431) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_430 | count_431)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_430 | idle_430) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_430 | idle_430)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_431 | count_432) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_431 | count_432)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_431 | idle_431) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_431 | idle_431)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_432 | count_433) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_432 | count_433)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_432 | idle_432) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_432 | idle_432)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_433 | count_434) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_433 | count_434)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_433 | idle_433) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_433 | idle_433)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_434 | count_435) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_434 | count_435)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_434 | idle_434) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_434 | idle_434)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_435 | count_436) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_435 | count_436)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_435 | idle_435) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_435 | idle_435)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_436 | count_437) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_436 | count_437)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_436 | idle_436) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_436 | idle_436)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_437 | count_438) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_437 | count_438)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_437 | idle_437) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_437 | idle_437)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_438 | count_439) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_438 | count_439)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_438 | idle_438) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_438 | idle_438)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_439 | count_440) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_439 | count_440)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_439 | idle_439) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_439 | idle_439)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_440 | count_441) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_440 | count_441)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_440 | idle_440) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_440 | idle_440)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_441 | count_442) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_441 | count_442)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_441 | idle_441) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_441 | idle_441)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_442 | count_443) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_442 | count_443)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_442 | idle_442) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_442 | idle_442)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_443 | count_444) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_443 | count_444)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_443 | idle_443) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_443 | idle_443)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_444 | count_445) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_444 | count_445)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_444 | idle_444) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_444 | idle_444)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_445 | count_446) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_445 | count_446)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_445 | idle_445) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_445 | idle_445)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_446 | count_447) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_446 | count_447)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_446 | idle_446) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_446 | idle_446)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_447 | count_448) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_447 | count_448)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_447 | idle_447) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_447 | idle_447)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_448 | count_449) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_448 | count_449)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_448 | idle_448) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_448 | idle_448)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_449 | count_450) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_449 | count_450)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_449 | idle_449) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_449 | idle_449)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_450 | count_451) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_450 | count_451)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_450 | idle_450) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_450 | idle_450)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_451 | count_452) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_451 | count_452)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_451 | idle_451) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_451 | idle_451)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_452 | count_453) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_452 | count_453)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_452 | idle_452) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_452 | idle_452)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_453 | count_454) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_453 | count_454)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_453 | idle_453) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_453 | idle_453)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_454 | count_455) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_454 | count_455)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_454 | idle_454) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_454 | idle_454)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_455 | count_456) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_455 | count_456)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_455 | idle_455) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_455 | idle_455)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_456 | count_457) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_456 | count_457)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_456 | idle_456) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_456 | idle_456)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_457 | count_458) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_457 | count_458)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_457 | idle_457) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_457 | idle_457)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_458 | count_459) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_458 | count_459)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_458 | idle_458) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_458 | idle_458)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_459 | count_460) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_459 | count_460)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_459 | idle_459) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_459 | idle_459)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_460 | count_461) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_460 | count_461)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_460 | idle_460) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_460 | idle_460)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_461 | count_462) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_461 | count_462)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_461 | idle_461) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_461 | idle_461)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_462 | count_463) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_462 | count_463)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_462 | idle_462) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_462 | idle_462)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_463 | count_464) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_463 | count_464)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_463 | idle_463) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_463 | idle_463)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_464 | count_465) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_464 | count_465)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_464 | idle_464) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_464 | idle_464)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_465 | count_466) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_465 | count_466)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_465 | idle_465) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_465 | idle_465)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_466 | count_467) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_466 | count_467)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_466 | idle_466) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_466 | idle_466)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_467 | count_468) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_467 | count_468)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_467 | idle_467) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_467 | idle_467)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_468 | count_469) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_468 | count_469)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_468 | idle_468) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_468 | idle_468)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_469 | count_470) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_469 | count_470)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_469 | idle_469) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_469 | idle_469)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_470 | count_471) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_470 | count_471)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_470 | idle_470) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_470 | idle_470)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_471 | count_472) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_471 | count_472)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_471 | idle_471) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_471 | idle_471)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_472 | count_473) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_472 | count_473)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_472 | idle_472) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_472 | idle_472)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_473 | count_474) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_473 | count_474)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_473 | idle_473) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_473 | idle_473)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_474 | count_475) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_474 | count_475)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_474 | idle_474) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_474 | idle_474)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_475 | count_476) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_475 | count_476)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_475 | idle_475) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_475 | idle_475)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_476 | count_477) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_476 | count_477)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_476 | idle_476) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_476 | idle_476)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_477 | count_478) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_477 | count_478)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_477 | idle_477) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_477 | idle_477)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_478 | count_479) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_478 | count_479)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_478 | idle_478) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_478 | idle_478)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_479 | count_480) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_479 | count_480)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_479 | idle_479) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_479 | idle_479)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_480 | count_481) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_480 | count_481)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_480 | idle_480) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_480 | idle_480)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_481 | count_482) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_481 | count_482)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_481 | idle_481) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_481 | idle_481)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_482 | count_483) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_482 | count_483)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_482 | idle_482) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_482 | idle_482)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_483 | count_484) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_483 | count_484)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_483 | idle_483) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_483 | idle_483)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_484 | count_485) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_484 | count_485)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_484 | idle_484) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_484 | idle_484)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_485 | count_486) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_485 | count_486)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_485 | idle_485) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_485 | idle_485)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_486 | count_487) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_486 | count_487)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_486 | idle_486) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_486 | idle_486)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_487 | count_488) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_487 | count_488)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_487 | idle_487) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_487 | idle_487)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_488 | count_489) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_488 | count_489)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_488 | idle_488) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_488 | idle_488)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_489 | count_490) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_489 | count_490)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_489 | idle_489) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_489 | idle_489)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_490 | count_491) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_490 | count_491)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_490 | idle_490) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_490 | idle_490)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_491 | count_492) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_491 | count_492)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_491 | idle_491) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_491 | idle_491)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_492 | count_493) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_492 | count_493)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_492 | idle_492) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_492 | idle_492)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_493 | count_494) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_493 | count_494)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_493 | idle_493) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_493 | idle_493)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_494 | count_495) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_494 | count_495)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_494 | idle_494) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_494 | idle_494)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_495 | count_496) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_495 | count_496)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_495 | idle_495) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_495 | idle_495)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_496 | count_497) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_496 | count_497)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_496 | idle_496) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_496 | idle_496)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_497 | count_498) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_497 | count_498)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_497 | idle_497) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_497 | idle_497)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_498 | count_499) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_498 | count_499)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_498 | idle_498) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_498 | idle_498)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_499 | count_500) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_499 | count_500)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_499 | idle_499) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_499 | idle_499)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_500 | count_501) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_500 | count_501)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_500 | idle_500) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_500 | idle_500)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_501 | count_502) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_501 | count_502)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_501 | idle_501) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_501 | idle_501)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_502 | count_503) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_502 | count_503)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_502 | idle_502) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_502 | idle_502)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_503 | count_504) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_503 | count_504)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_503 | idle_503) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_503 | idle_503)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_504 | count_505) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_504 | count_505)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_504 | idle_504) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_504 | idle_504)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_505 | count_506) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_505 | count_506)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_505 | idle_505) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_505 | idle_505)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_506 | count_507) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_506 | count_507)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_506 | idle_506) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_506 | idle_506)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_507 | count_508) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_507 | count_508)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_507 | idle_507) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_507 | idle_507)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_508 | count_509) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_508 | count_509)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_508 | idle_508) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_508 | idle_508)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_509 | count_510) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_509 | count_510)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_509 | idle_509) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_509 | idle_509)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_510 | count_511) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_510 | count_511)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_510 | idle_510) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_510 | idle_510)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~dec_511 | count_512) & ~reset) begin
          $fatal; // @[ToAXI4.scala 262:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_511 | count_512)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:262 assert (!dec || count =/= UInt(0))        // underflow\n"); // @[ToAXI4.scala 262:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~inc_511 | idle_511) & _T_10) begin
          $fatal; // @[ToAXI4.scala 263:16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_511 | idle_511)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:263 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); // @[ToAXI4.scala 263:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    TLToAXI4_covState <= TLToAXI4_xor0;
    if (TLToAXI4_covMap_write_en & TLToAXI4_covMap_write_mask) begin
      TLToAXI4_covMap[TLToAXI4_covMap_write_addr] <= TLToAXI4_covMap_write_data; // @[Coverage map for TLToAXI4]
    end
    if (!(TLToAXI4_covMap_read_data | metaReset)) begin
      TLToAXI4_covSum <= TLToAXI4_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_519 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    TLToAXI4_covMap[initvar] = 0; //_519[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count_512 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  count_511 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  count_510 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  count_509 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  count_508 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  count_507 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  count_506 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  count_505 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  count_504 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  count_503 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  count_502 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  count_501 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  count_500 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  count_499 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  count_498 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  count_497 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  count_496 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  count_495 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  count_494 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  count_493 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  count_492 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  count_491 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  count_490 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  count_489 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  count_488 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  count_487 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  count_486 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  count_485 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  count_484 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  count_483 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  count_482 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  count_481 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  count_480 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  count_479 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  count_478 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  count_477 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  count_476 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  count_475 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  count_474 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  count_473 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  count_472 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  count_471 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  count_470 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  count_469 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  count_468 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  count_467 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  count_466 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  count_465 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  count_464 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  count_463 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  count_462 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  count_461 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  count_460 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  count_459 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  count_458 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  count_457 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  count_456 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  count_455 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  count_454 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  count_453 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  count_452 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  count_451 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  count_450 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  count_449 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  count_448 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  count_447 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  count_446 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  count_445 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  count_444 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  count_443 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  count_442 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  count_441 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  count_440 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  count_439 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  count_438 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  count_437 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  count_436 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  count_435 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  count_434 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  count_433 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  count_432 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  count_431 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  count_430 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  count_429 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  count_428 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  count_427 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  count_426 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  count_425 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  count_424 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  count_423 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  count_422 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  count_421 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  count_420 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  count_419 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  count_418 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  count_417 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  count_416 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  count_415 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  count_414 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  count_413 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  count_412 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  count_411 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  count_410 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  count_409 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  count_408 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  count_407 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  count_406 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  count_405 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  count_404 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  count_403 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  count_402 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  count_401 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  count_400 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  count_399 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  count_398 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  count_397 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  count_396 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  count_395 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  count_394 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  count_393 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  count_392 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  count_391 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  count_390 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  count_389 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  count_388 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  count_387 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  count_386 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  count_385 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  count_384 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  count_383 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  count_382 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  count_381 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  count_380 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  count_379 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  count_378 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  count_377 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  count_376 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  count_375 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  count_374 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  count_373 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  count_372 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  count_371 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  count_370 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  count_369 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  count_368 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  count_367 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  count_366 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  count_365 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  count_364 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  count_363 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  count_362 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  count_361 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  count_360 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  count_359 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  count_358 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  count_357 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  count_356 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  count_355 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  count_354 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  count_353 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  count_352 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  count_351 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  count_350 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  count_349 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  count_348 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  count_347 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  count_346 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  count_345 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  count_344 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  count_343 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  count_342 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  count_341 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  count_340 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  count_339 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  count_338 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  count_337 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  count_336 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  count_335 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  count_334 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  count_333 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  count_332 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  count_331 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  count_330 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  count_329 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  count_328 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  count_327 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  count_326 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  count_325 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  count_324 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  count_323 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  count_322 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  count_321 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  count_320 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  count_319 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  count_318 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  count_317 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  count_316 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  count_315 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  count_314 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  count_313 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  count_312 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  count_311 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  count_310 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  count_309 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  count_308 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  count_307 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  count_306 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  count_305 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  count_304 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  count_303 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  count_302 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  count_301 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  count_300 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  count_299 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  count_298 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  count_297 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  count_296 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  count_295 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  count_294 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  count_293 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  count_292 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  count_291 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  count_290 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  count_289 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  count_288 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  count_287 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  count_286 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  count_285 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  count_284 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  count_283 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  count_282 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  count_281 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  count_280 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  count_279 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  count_278 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  count_277 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  count_276 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  count_275 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  count_274 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  count_273 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  count_272 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  count_271 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  count_270 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  count_269 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  count_268 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  count_267 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  count_266 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  count_265 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  count_264 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  count_263 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  count_262 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  count_261 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  count_260 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  count_259 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  count_258 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  count_257 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  count_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  count_255 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  count_254 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  count_253 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  count_252 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  count_251 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  count_250 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  count_249 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  count_248 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  count_247 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  count_246 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  count_245 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  count_244 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  count_243 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  count_242 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  count_241 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  count_240 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  count_239 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  count_238 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  count_237 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  count_236 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  count_235 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  count_234 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  count_233 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  count_232 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  count_231 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  count_230 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  count_229 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  count_228 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  count_227 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  count_226 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  count_225 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  count_224 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  count_223 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  count_222 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  count_221 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  count_220 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  count_219 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  count_218 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  count_217 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  count_216 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  count_215 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  count_214 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  count_213 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  count_212 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  count_211 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  count_210 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  count_209 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  count_208 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  count_207 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  count_206 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  count_205 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  count_204 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  count_203 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  count_202 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  count_201 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  count_200 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  count_199 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  count_198 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  count_197 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  count_196 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  count_195 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  count_194 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  count_193 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  count_192 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  count_191 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  count_190 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  count_189 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  count_188 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  count_187 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  count_186 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  count_185 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  count_184 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  count_183 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  count_182 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  count_181 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  count_180 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  count_179 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  count_178 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  count_177 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  count_176 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  count_175 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  count_174 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  count_173 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  count_172 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  count_171 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  count_170 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  count_169 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  count_168 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  count_167 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  count_166 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  count_165 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  count_164 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  count_163 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  count_162 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  count_161 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  count_160 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  count_159 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  count_158 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  count_157 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  count_156 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  count_155 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  count_154 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  count_153 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  count_152 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  count_151 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  count_150 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  count_149 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  count_148 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  count_147 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  count_146 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  count_145 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  count_144 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  count_143 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  count_142 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  count_141 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  count_140 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  count_139 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  count_138 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  count_137 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  count_136 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  count_135 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  count_134 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  count_133 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  count_132 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  count_131 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  count_130 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  count_129 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  count_128 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  count_127 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  count_126 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  count_125 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  count_124 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  count_123 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  count_122 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  count_121 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  count_120 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  count_119 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  count_118 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  count_117 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  count_116 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  count_115 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  count_114 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  count_113 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  count_112 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  count_111 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  count_110 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  count_109 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  count_108 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  count_107 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  count_106 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  count_105 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  count_104 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  count_103 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  count_102 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  count_101 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  count_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  count_99 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  count_98 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  count_97 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  count_96 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  count_95 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  count_94 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  count_93 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  count_92 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  count_91 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  count_90 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  count_89 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  count_88 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  count_87 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  count_86 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  count_85 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  count_84 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  count_83 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  count_82 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  count_81 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  count_80 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  count_79 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  count_78 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  count_77 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  count_76 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  count_75 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  count_74 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  count_73 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  count_72 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  count_71 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  count_70 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  count_69 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  count_68 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  count_67 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  count_66 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  count_65 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  count_64 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  count_63 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  count_62 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  count_61 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  count_60 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  count_59 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  count_58 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  count_57 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  count_56 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  count_55 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  count_54 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  count_53 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  count_52 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  count_51 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  count_50 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  count_49 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  count_48 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  count_47 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  count_46 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  count_45 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  count_44 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  count_43 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  count_42 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  count_41 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  count_40 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  count_39 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  count_38 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  count_37 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  count_36 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  count_35 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  count_34 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  count_33 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  count_32 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  count_31 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  count_30 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  count_29 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  count_28 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  count_27 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  count_26 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  count_25 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  count_24 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  count_23 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  count_22 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  count_21 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  count_20 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  count_19 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  count_18 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  count_17 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  count_16 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  count_15 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  count_14 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  count_13 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  count_12 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  count_11 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  count_10 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  count_9 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  count_8 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  count_7 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  count_6 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  count_5 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  count_4 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  count_3 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  count_2 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  count_1 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  counter = _RAND_512[2:0];
  _RAND_513 = {1{`RANDOM}};
  doneAW = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  r_holds_d = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  b_delay = _RAND_515[2:0];
  _RAND_516 = {1{`RANDOM}};
  r_first = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  r_denied_r = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  TLToAXI4_covState = 0; //_518[19:0];
  _RAND_520 = {1{`RANDOM}};
  TLToAXI4_covSum = 0; //_520[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLInterconnectCoupler_13(
  input         clock,
  input         reset,
  input         auto_axi4yank_out_aw_ready,
  output        auto_axi4yank_out_aw_valid,
  output [3:0]  auto_axi4yank_out_aw_bits_id,
  output [31:0] auto_axi4yank_out_aw_bits_addr,
  output [7:0]  auto_axi4yank_out_aw_bits_len,
  output [2:0]  auto_axi4yank_out_aw_bits_size,
  output [1:0]  auto_axi4yank_out_aw_bits_burst,
  output        auto_axi4yank_out_aw_bits_lock,
  output [3:0]  auto_axi4yank_out_aw_bits_cache,
  output [2:0]  auto_axi4yank_out_aw_bits_prot,
  output [3:0]  auto_axi4yank_out_aw_bits_qos,
  input         auto_axi4yank_out_w_ready,
  output        auto_axi4yank_out_w_valid,
  output [63:0] auto_axi4yank_out_w_bits_data,
  output [7:0]  auto_axi4yank_out_w_bits_strb,
  output        auto_axi4yank_out_w_bits_last,
  output        auto_axi4yank_out_b_ready,
  input         auto_axi4yank_out_b_valid,
  input  [3:0]  auto_axi4yank_out_b_bits_id,
  input  [1:0]  auto_axi4yank_out_b_bits_resp,
  input         auto_axi4yank_out_ar_ready,
  output        auto_axi4yank_out_ar_valid,
  output [3:0]  auto_axi4yank_out_ar_bits_id,
  output [31:0] auto_axi4yank_out_ar_bits_addr,
  output [7:0]  auto_axi4yank_out_ar_bits_len,
  output [2:0]  auto_axi4yank_out_ar_bits_size,
  output [1:0]  auto_axi4yank_out_ar_bits_burst,
  output        auto_axi4yank_out_ar_bits_lock,
  output [3:0]  auto_axi4yank_out_ar_bits_cache,
  output [2:0]  auto_axi4yank_out_ar_bits_prot,
  output [3:0]  auto_axi4yank_out_ar_bits_qos,
  output        auto_axi4yank_out_r_ready,
  input         auto_axi4yank_out_r_valid,
  input  [3:0]  auto_axi4yank_out_r_bits_id,
  input  [63:0] auto_axi4yank_out_r_bits_data,
  input  [1:0]  auto_axi4yank_out_r_bits_resp,
  input         auto_axi4yank_out_r_bits_last,
  output        auto_tl_in_a_ready,
  input         auto_tl_in_a_valid,
  input  [2:0]  auto_tl_in_a_bits_opcode,
  input  [2:0]  auto_tl_in_a_bits_size,
  input  [8:0]  auto_tl_in_a_bits_source,
  input  [31:0] auto_tl_in_a_bits_address,
  input         auto_tl_in_a_bits_user_amba_prot_bufferable,
  input         auto_tl_in_a_bits_user_amba_prot_modifiable,
  input         auto_tl_in_a_bits_user_amba_prot_readalloc,
  input         auto_tl_in_a_bits_user_amba_prot_writealloc,
  input         auto_tl_in_a_bits_user_amba_prot_privileged,
  input         auto_tl_in_a_bits_user_amba_prot_secure,
  input         auto_tl_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_tl_in_a_bits_mask,
  input  [63:0] auto_tl_in_a_bits_data,
  input         auto_tl_in_d_ready,
  output        auto_tl_in_d_valid,
  output [2:0]  auto_tl_in_d_bits_opcode,
  output [2:0]  auto_tl_in_d_bits_size,
  output [8:0]  auto_tl_in_d_bits_source,
  output        auto_tl_in_d_bits_denied,
  output [63:0] auto_tl_in_d_bits_data,
  output        auto_tl_in_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  axi4yank_clock; // @[UserYanker.scala 105:30]
  wire  axi4yank_reset; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_aw_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_in_aw_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_aw_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_aw_bits_size; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_aw_bits_burst; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_bits_lock; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_aw_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_aw_bits_prot; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_aw_bits_qos; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_aw_bits_echo_tl_state_size; // @[UserYanker.scala 105:30]
  wire [8:0] axi4yank_auto_in_aw_bits_echo_tl_state_source; // @[UserYanker.scala 105:30]
  wire [4:0] axi4yank_auto_in_aw_bits_echo_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_w_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_w_valid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_in_w_bits_data; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_w_bits_strb; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_w_bits_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_b_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_b_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_b_bits_id; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_b_bits_resp; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_b_bits_echo_tl_state_size; // @[UserYanker.scala 105:30]
  wire [8:0] axi4yank_auto_in_b_bits_echo_tl_state_source; // @[UserYanker.scala 105:30]
  wire [4:0] axi4yank_auto_in_b_bits_echo_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_ar_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_in_ar_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_ar_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_ar_bits_size; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_ar_bits_burst; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_bits_lock; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_ar_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_ar_bits_prot; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_ar_bits_qos; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_ar_bits_echo_tl_state_size; // @[UserYanker.scala 105:30]
  wire [8:0] axi4yank_auto_in_ar_bits_echo_tl_state_source; // @[UserYanker.scala 105:30]
  wire [4:0] axi4yank_auto_in_ar_bits_echo_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_r_bits_id; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_in_r_bits_data; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_r_bits_resp; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_r_bits_echo_tl_state_size; // @[UserYanker.scala 105:30]
  wire [8:0] axi4yank_auto_in_r_bits_echo_tl_state_source; // @[UserYanker.scala 105:30]
  wire [4:0] axi4yank_auto_in_r_bits_echo_extra_id; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_bits_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_aw_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_aw_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_aw_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_out_aw_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_aw_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_aw_bits_size; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_aw_bits_burst; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_aw_bits_lock; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_aw_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_aw_bits_prot; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_aw_bits_qos; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_w_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_w_valid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_out_w_bits_data; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_w_bits_strb; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_w_bits_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_b_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_b_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_b_bits_id; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_b_bits_resp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_ar_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_ar_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_ar_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_out_ar_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_ar_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_ar_bits_size; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_ar_bits_burst; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_ar_bits_lock; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_ar_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_ar_bits_prot; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_ar_bits_qos; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_r_bits_id; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_out_r_bits_data; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_r_bits_resp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_bits_last; // @[UserYanker.scala 105:30]
  wire [29:0] axi4yank_io_covSum; // @[UserYanker.scala 105:30]
  wire  axi4index_auto_in_aw_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_aw_valid; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_in_aw_bits_id; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_in_aw_bits_addr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_aw_bits_len; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_aw_bits_size; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_aw_bits_burst; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_aw_bits_lock; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_aw_bits_cache; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_aw_bits_prot; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_aw_bits_qos; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_aw_bits_echo_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_in_aw_bits_echo_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_w_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_w_valid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_in_w_bits_data; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_w_bits_strb; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_w_bits_last; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_b_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_b_valid; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_in_b_bits_id; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_b_bits_resp; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_b_bits_echo_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_in_b_bits_echo_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_ar_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_ar_valid; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_in_ar_bits_id; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_in_ar_bits_addr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_in_ar_bits_len; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_ar_bits_size; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_ar_bits_burst; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_ar_bits_lock; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_ar_bits_cache; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_in_ar_bits_prot; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_ar_bits_qos; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_ar_bits_echo_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_in_ar_bits_echo_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_r_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_r_valid; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_in_r_bits_id; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_in_r_bits_data; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_in_r_bits_resp; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_in_r_bits_echo_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_in_r_bits_echo_tl_state_source; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_in_r_bits_last; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_aw_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_aw_valid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_aw_bits_id; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_out_aw_bits_addr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_out_aw_bits_len; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_aw_bits_size; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_aw_bits_burst; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_aw_bits_lock; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_aw_bits_cache; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_aw_bits_prot; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_aw_bits_qos; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_aw_bits_echo_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_out_aw_bits_echo_tl_state_source; // @[IdIndexer.scala 91:31]
  wire [4:0] axi4index_auto_out_aw_bits_echo_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_w_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_w_valid; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_out_w_bits_data; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_out_w_bits_strb; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_w_bits_last; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_b_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_b_valid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_b_bits_id; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_b_bits_resp; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_b_bits_echo_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_out_b_bits_echo_tl_state_source; // @[IdIndexer.scala 91:31]
  wire [4:0] axi4index_auto_out_b_bits_echo_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_ar_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_ar_valid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_ar_bits_id; // @[IdIndexer.scala 91:31]
  wire [31:0] axi4index_auto_out_ar_bits_addr; // @[IdIndexer.scala 91:31]
  wire [7:0] axi4index_auto_out_ar_bits_len; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_ar_bits_size; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_ar_bits_burst; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_ar_bits_lock; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_ar_bits_cache; // @[IdIndexer.scala 91:31]
  wire [2:0] axi4index_auto_out_ar_bits_prot; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_ar_bits_qos; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_ar_bits_echo_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_out_ar_bits_echo_tl_state_source; // @[IdIndexer.scala 91:31]
  wire [4:0] axi4index_auto_out_ar_bits_echo_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_r_ready; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_r_valid; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_r_bits_id; // @[IdIndexer.scala 91:31]
  wire [63:0] axi4index_auto_out_r_bits_data; // @[IdIndexer.scala 91:31]
  wire [1:0] axi4index_auto_out_r_bits_resp; // @[IdIndexer.scala 91:31]
  wire [3:0] axi4index_auto_out_r_bits_echo_tl_state_size; // @[IdIndexer.scala 91:31]
  wire [8:0] axi4index_auto_out_r_bits_echo_tl_state_source; // @[IdIndexer.scala 91:31]
  wire [4:0] axi4index_auto_out_r_bits_echo_extra_id; // @[IdIndexer.scala 91:31]
  wire  axi4index_auto_out_r_bits_last; // @[IdIndexer.scala 91:31]
  wire [29:0] axi4index_io_covSum; // @[IdIndexer.scala 91:31]
  wire  tl2axi4_clock; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_reset; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_ready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_valid; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_in_a_bits_opcode; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_in_a_bits_size; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_in_a_bits_source; // @[ToAXI4.scala 283:29]
  wire [31:0] tl2axi4_auto_in_a_bits_address; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_bits_user_amba_prot_bufferable; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_bits_user_amba_prot_modifiable; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_bits_user_amba_prot_readalloc; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_bits_user_amba_prot_writealloc; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_bits_user_amba_prot_privileged; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_bits_user_amba_prot_secure; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_a_bits_user_amba_prot_fetch; // @[ToAXI4.scala 283:29]
  wire [7:0] tl2axi4_auto_in_a_bits_mask; // @[ToAXI4.scala 283:29]
  wire [63:0] tl2axi4_auto_in_a_bits_data; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_d_ready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_d_valid; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_in_d_bits_opcode; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_in_d_bits_size; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_in_d_bits_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_d_bits_denied; // @[ToAXI4.scala 283:29]
  wire [63:0] tl2axi4_auto_in_d_bits_data; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_in_d_bits_corrupt; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_aw_ready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_aw_valid; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_out_aw_bits_id; // @[ToAXI4.scala 283:29]
  wire [31:0] tl2axi4_auto_out_aw_bits_addr; // @[ToAXI4.scala 283:29]
  wire [7:0] tl2axi4_auto_out_aw_bits_len; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_out_aw_bits_size; // @[ToAXI4.scala 283:29]
  wire [1:0] tl2axi4_auto_out_aw_bits_burst; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_aw_bits_lock; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_aw_bits_cache; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_out_aw_bits_prot; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_aw_bits_qos; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_aw_bits_echo_tl_state_size; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_out_aw_bits_echo_tl_state_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_w_ready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_w_valid; // @[ToAXI4.scala 283:29]
  wire [63:0] tl2axi4_auto_out_w_bits_data; // @[ToAXI4.scala 283:29]
  wire [7:0] tl2axi4_auto_out_w_bits_strb; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_w_bits_last; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_b_ready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_b_valid; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_out_b_bits_id; // @[ToAXI4.scala 283:29]
  wire [1:0] tl2axi4_auto_out_b_bits_resp; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_b_bits_echo_tl_state_size; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_out_b_bits_echo_tl_state_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_ar_ready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_ar_valid; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_out_ar_bits_id; // @[ToAXI4.scala 283:29]
  wire [31:0] tl2axi4_auto_out_ar_bits_addr; // @[ToAXI4.scala 283:29]
  wire [7:0] tl2axi4_auto_out_ar_bits_len; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_out_ar_bits_size; // @[ToAXI4.scala 283:29]
  wire [1:0] tl2axi4_auto_out_ar_bits_burst; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_ar_bits_lock; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_ar_bits_cache; // @[ToAXI4.scala 283:29]
  wire [2:0] tl2axi4_auto_out_ar_bits_prot; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_ar_bits_qos; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_ar_bits_echo_tl_state_size; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_out_ar_bits_echo_tl_state_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_r_ready; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_r_valid; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_out_r_bits_id; // @[ToAXI4.scala 283:29]
  wire [63:0] tl2axi4_auto_out_r_bits_data; // @[ToAXI4.scala 283:29]
  wire [1:0] tl2axi4_auto_out_r_bits_resp; // @[ToAXI4.scala 283:29]
  wire [3:0] tl2axi4_auto_out_r_bits_echo_tl_state_size; // @[ToAXI4.scala 283:29]
  wire [8:0] tl2axi4_auto_out_r_bits_echo_tl_state_source; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_auto_out_r_bits_last; // @[ToAXI4.scala 283:29]
  wire [29:0] tl2axi4_io_covSum; // @[ToAXI4.scala 283:29]
  wire  tl2axi4_metaReset; // @[ToAXI4.scala 283:29]
  wire  widget_auto_in_a_ready;
  wire  widget_auto_in_a_valid;
  wire [2:0] widget_auto_in_a_bits_opcode;
  wire [2:0] widget_auto_in_a_bits_size;
  wire [8:0] widget_auto_in_a_bits_source;
  wire [31:0] widget_auto_in_a_bits_address;
  wire  widget_auto_in_a_bits_user_amba_prot_bufferable;
  wire  widget_auto_in_a_bits_user_amba_prot_modifiable;
  wire  widget_auto_in_a_bits_user_amba_prot_readalloc;
  wire  widget_auto_in_a_bits_user_amba_prot_writealloc;
  wire  widget_auto_in_a_bits_user_amba_prot_privileged;
  wire  widget_auto_in_a_bits_user_amba_prot_secure;
  wire  widget_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] widget_auto_in_a_bits_mask;
  wire [63:0] widget_auto_in_a_bits_data;
  wire  widget_auto_in_d_ready;
  wire  widget_auto_in_d_valid;
  wire [2:0] widget_auto_in_d_bits_opcode;
  wire [2:0] widget_auto_in_d_bits_size;
  wire [8:0] widget_auto_in_d_bits_source;
  wire  widget_auto_in_d_bits_denied;
  wire [63:0] widget_auto_in_d_bits_data;
  wire  widget_auto_in_d_bits_corrupt;
  wire  widget_auto_out_a_ready;
  wire  widget_auto_out_a_valid;
  wire [2:0] widget_auto_out_a_bits_opcode;
  wire [2:0] widget_auto_out_a_bits_size;
  wire [8:0] widget_auto_out_a_bits_source;
  wire [31:0] widget_auto_out_a_bits_address;
  wire  widget_auto_out_a_bits_user_amba_prot_bufferable;
  wire  widget_auto_out_a_bits_user_amba_prot_modifiable;
  wire  widget_auto_out_a_bits_user_amba_prot_readalloc;
  wire  widget_auto_out_a_bits_user_amba_prot_writealloc;
  wire  widget_auto_out_a_bits_user_amba_prot_privileged;
  wire  widget_auto_out_a_bits_user_amba_prot_secure;
  wire  widget_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] widget_auto_out_a_bits_mask;
  wire [63:0] widget_auto_out_a_bits_data;
  wire  widget_auto_out_d_ready;
  wire  widget_auto_out_d_valid;
  wire [2:0] widget_auto_out_d_bits_opcode;
  wire [2:0] widget_auto_out_d_bits_size;
  wire [8:0] widget_auto_out_d_bits_source;
  wire  widget_auto_out_d_bits_denied;
  wire [63:0] widget_auto_out_d_bits_data;
  wire  widget_auto_out_d_bits_corrupt;
  wire [29:0] TLInterconnectCoupler_13_covSum;
  wire [29:0] axi4yank_sum;
  wire [29:0] axi4index_sum;
  wire [29:0] tl2axi4_sum;
  AXI4UserYanker_1 axi4yank ( // @[UserYanker.scala 105:30]
    .clock(axi4yank_clock),
    .reset(axi4yank_reset),
    .auto_in_aw_ready(axi4yank_auto_in_aw_ready),
    .auto_in_aw_valid(axi4yank_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4yank_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4yank_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4yank_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4yank_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4yank_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4yank_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4yank_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4yank_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4yank_auto_in_aw_bits_qos),
    .auto_in_aw_bits_echo_tl_state_size(axi4yank_auto_in_aw_bits_echo_tl_state_size),
    .auto_in_aw_bits_echo_tl_state_source(axi4yank_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_aw_bits_echo_extra_id(axi4yank_auto_in_aw_bits_echo_extra_id),
    .auto_in_w_ready(axi4yank_auto_in_w_ready),
    .auto_in_w_valid(axi4yank_auto_in_w_valid),
    .auto_in_w_bits_data(axi4yank_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4yank_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4yank_auto_in_w_bits_last),
    .auto_in_b_ready(axi4yank_auto_in_b_ready),
    .auto_in_b_valid(axi4yank_auto_in_b_valid),
    .auto_in_b_bits_id(axi4yank_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4yank_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_tl_state_size(axi4yank_auto_in_b_bits_echo_tl_state_size),
    .auto_in_b_bits_echo_tl_state_source(axi4yank_auto_in_b_bits_echo_tl_state_source),
    .auto_in_b_bits_echo_extra_id(axi4yank_auto_in_b_bits_echo_extra_id),
    .auto_in_ar_ready(axi4yank_auto_in_ar_ready),
    .auto_in_ar_valid(axi4yank_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4yank_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4yank_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4yank_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4yank_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4yank_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4yank_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4yank_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4yank_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4yank_auto_in_ar_bits_qos),
    .auto_in_ar_bits_echo_tl_state_size(axi4yank_auto_in_ar_bits_echo_tl_state_size),
    .auto_in_ar_bits_echo_tl_state_source(axi4yank_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_ar_bits_echo_extra_id(axi4yank_auto_in_ar_bits_echo_extra_id),
    .auto_in_r_ready(axi4yank_auto_in_r_ready),
    .auto_in_r_valid(axi4yank_auto_in_r_valid),
    .auto_in_r_bits_id(axi4yank_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4yank_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4yank_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_tl_state_size(axi4yank_auto_in_r_bits_echo_tl_state_size),
    .auto_in_r_bits_echo_tl_state_source(axi4yank_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_echo_extra_id(axi4yank_auto_in_r_bits_echo_extra_id),
    .auto_in_r_bits_last(axi4yank_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4yank_auto_out_aw_ready),
    .auto_out_aw_valid(axi4yank_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4yank_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4yank_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4yank_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4yank_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4yank_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4yank_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4yank_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4yank_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4yank_auto_out_aw_bits_qos),
    .auto_out_w_ready(axi4yank_auto_out_w_ready),
    .auto_out_w_valid(axi4yank_auto_out_w_valid),
    .auto_out_w_bits_data(axi4yank_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4yank_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4yank_auto_out_w_bits_last),
    .auto_out_b_ready(axi4yank_auto_out_b_ready),
    .auto_out_b_valid(axi4yank_auto_out_b_valid),
    .auto_out_b_bits_id(axi4yank_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4yank_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4yank_auto_out_ar_ready),
    .auto_out_ar_valid(axi4yank_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4yank_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4yank_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4yank_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4yank_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4yank_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4yank_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4yank_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4yank_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4yank_auto_out_ar_bits_qos),
    .auto_out_r_ready(axi4yank_auto_out_r_ready),
    .auto_out_r_valid(axi4yank_auto_out_r_valid),
    .auto_out_r_bits_id(axi4yank_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4yank_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4yank_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4yank_auto_out_r_bits_last),
    .io_covSum(axi4yank_io_covSum)
  );
  AXI4IdIndexer_1 axi4index ( // @[IdIndexer.scala 91:31]
    .auto_in_aw_ready(axi4index_auto_in_aw_ready),
    .auto_in_aw_valid(axi4index_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4index_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4index_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4index_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4index_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4index_auto_in_aw_bits_burst),
    .auto_in_aw_bits_lock(axi4index_auto_in_aw_bits_lock),
    .auto_in_aw_bits_cache(axi4index_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4index_auto_in_aw_bits_prot),
    .auto_in_aw_bits_qos(axi4index_auto_in_aw_bits_qos),
    .auto_in_aw_bits_echo_tl_state_size(axi4index_auto_in_aw_bits_echo_tl_state_size),
    .auto_in_aw_bits_echo_tl_state_source(axi4index_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_w_ready(axi4index_auto_in_w_ready),
    .auto_in_w_valid(axi4index_auto_in_w_valid),
    .auto_in_w_bits_data(axi4index_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4index_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4index_auto_in_w_bits_last),
    .auto_in_b_ready(axi4index_auto_in_b_ready),
    .auto_in_b_valid(axi4index_auto_in_b_valid),
    .auto_in_b_bits_id(axi4index_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4index_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_tl_state_size(axi4index_auto_in_b_bits_echo_tl_state_size),
    .auto_in_b_bits_echo_tl_state_source(axi4index_auto_in_b_bits_echo_tl_state_source),
    .auto_in_ar_ready(axi4index_auto_in_ar_ready),
    .auto_in_ar_valid(axi4index_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4index_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4index_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4index_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4index_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4index_auto_in_ar_bits_burst),
    .auto_in_ar_bits_lock(axi4index_auto_in_ar_bits_lock),
    .auto_in_ar_bits_cache(axi4index_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4index_auto_in_ar_bits_prot),
    .auto_in_ar_bits_qos(axi4index_auto_in_ar_bits_qos),
    .auto_in_ar_bits_echo_tl_state_size(axi4index_auto_in_ar_bits_echo_tl_state_size),
    .auto_in_ar_bits_echo_tl_state_source(axi4index_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_r_ready(axi4index_auto_in_r_ready),
    .auto_in_r_valid(axi4index_auto_in_r_valid),
    .auto_in_r_bits_id(axi4index_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4index_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4index_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_tl_state_size(axi4index_auto_in_r_bits_echo_tl_state_size),
    .auto_in_r_bits_echo_tl_state_source(axi4index_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_last(axi4index_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4index_auto_out_aw_ready),
    .auto_out_aw_valid(axi4index_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4index_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4index_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4index_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4index_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4index_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(axi4index_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(axi4index_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4index_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(axi4index_auto_out_aw_bits_qos),
    .auto_out_aw_bits_echo_tl_state_size(axi4index_auto_out_aw_bits_echo_tl_state_size),
    .auto_out_aw_bits_echo_tl_state_source(axi4index_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_aw_bits_echo_extra_id(axi4index_auto_out_aw_bits_echo_extra_id),
    .auto_out_w_ready(axi4index_auto_out_w_ready),
    .auto_out_w_valid(axi4index_auto_out_w_valid),
    .auto_out_w_bits_data(axi4index_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4index_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4index_auto_out_w_bits_last),
    .auto_out_b_ready(axi4index_auto_out_b_ready),
    .auto_out_b_valid(axi4index_auto_out_b_valid),
    .auto_out_b_bits_id(axi4index_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4index_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_tl_state_size(axi4index_auto_out_b_bits_echo_tl_state_size),
    .auto_out_b_bits_echo_tl_state_source(axi4index_auto_out_b_bits_echo_tl_state_source),
    .auto_out_b_bits_echo_extra_id(axi4index_auto_out_b_bits_echo_extra_id),
    .auto_out_ar_ready(axi4index_auto_out_ar_ready),
    .auto_out_ar_valid(axi4index_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4index_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4index_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4index_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4index_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4index_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(axi4index_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(axi4index_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4index_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(axi4index_auto_out_ar_bits_qos),
    .auto_out_ar_bits_echo_tl_state_size(axi4index_auto_out_ar_bits_echo_tl_state_size),
    .auto_out_ar_bits_echo_tl_state_source(axi4index_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_ar_bits_echo_extra_id(axi4index_auto_out_ar_bits_echo_extra_id),
    .auto_out_r_ready(axi4index_auto_out_r_ready),
    .auto_out_r_valid(axi4index_auto_out_r_valid),
    .auto_out_r_bits_id(axi4index_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4index_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4index_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_tl_state_size(axi4index_auto_out_r_bits_echo_tl_state_size),
    .auto_out_r_bits_echo_tl_state_source(axi4index_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_echo_extra_id(axi4index_auto_out_r_bits_echo_extra_id),
    .auto_out_r_bits_last(axi4index_auto_out_r_bits_last),
    .io_covSum(axi4index_io_covSum)
  );
  TLToAXI4 tl2axi4 ( // @[ToAXI4.scala 283:29]
    .clock(tl2axi4_clock),
    .reset(tl2axi4_reset),
    .auto_in_a_ready(tl2axi4_auto_in_a_ready),
    .auto_in_a_valid(tl2axi4_auto_in_a_valid),
    .auto_in_a_bits_opcode(tl2axi4_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(tl2axi4_auto_in_a_bits_size),
    .auto_in_a_bits_source(tl2axi4_auto_in_a_bits_source),
    .auto_in_a_bits_address(tl2axi4_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(tl2axi4_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(tl2axi4_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(tl2axi4_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(tl2axi4_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(tl2axi4_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(tl2axi4_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(tl2axi4_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(tl2axi4_auto_in_a_bits_mask),
    .auto_in_a_bits_data(tl2axi4_auto_in_a_bits_data),
    .auto_in_d_ready(tl2axi4_auto_in_d_ready),
    .auto_in_d_valid(tl2axi4_auto_in_d_valid),
    .auto_in_d_bits_opcode(tl2axi4_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(tl2axi4_auto_in_d_bits_size),
    .auto_in_d_bits_source(tl2axi4_auto_in_d_bits_source),
    .auto_in_d_bits_denied(tl2axi4_auto_in_d_bits_denied),
    .auto_in_d_bits_data(tl2axi4_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(tl2axi4_auto_in_d_bits_corrupt),
    .auto_out_aw_ready(tl2axi4_auto_out_aw_ready),
    .auto_out_aw_valid(tl2axi4_auto_out_aw_valid),
    .auto_out_aw_bits_id(tl2axi4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(tl2axi4_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(tl2axi4_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(tl2axi4_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(tl2axi4_auto_out_aw_bits_burst),
    .auto_out_aw_bits_lock(tl2axi4_auto_out_aw_bits_lock),
    .auto_out_aw_bits_cache(tl2axi4_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(tl2axi4_auto_out_aw_bits_prot),
    .auto_out_aw_bits_qos(tl2axi4_auto_out_aw_bits_qos),
    .auto_out_aw_bits_echo_tl_state_size(tl2axi4_auto_out_aw_bits_echo_tl_state_size),
    .auto_out_aw_bits_echo_tl_state_source(tl2axi4_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_w_ready(tl2axi4_auto_out_w_ready),
    .auto_out_w_valid(tl2axi4_auto_out_w_valid),
    .auto_out_w_bits_data(tl2axi4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(tl2axi4_auto_out_w_bits_strb),
    .auto_out_w_bits_last(tl2axi4_auto_out_w_bits_last),
    .auto_out_b_ready(tl2axi4_auto_out_b_ready),
    .auto_out_b_valid(tl2axi4_auto_out_b_valid),
    .auto_out_b_bits_id(tl2axi4_auto_out_b_bits_id),
    .auto_out_b_bits_resp(tl2axi4_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_tl_state_size(tl2axi4_auto_out_b_bits_echo_tl_state_size),
    .auto_out_b_bits_echo_tl_state_source(tl2axi4_auto_out_b_bits_echo_tl_state_source),
    .auto_out_ar_ready(tl2axi4_auto_out_ar_ready),
    .auto_out_ar_valid(tl2axi4_auto_out_ar_valid),
    .auto_out_ar_bits_id(tl2axi4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(tl2axi4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(tl2axi4_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(tl2axi4_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(tl2axi4_auto_out_ar_bits_burst),
    .auto_out_ar_bits_lock(tl2axi4_auto_out_ar_bits_lock),
    .auto_out_ar_bits_cache(tl2axi4_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(tl2axi4_auto_out_ar_bits_prot),
    .auto_out_ar_bits_qos(tl2axi4_auto_out_ar_bits_qos),
    .auto_out_ar_bits_echo_tl_state_size(tl2axi4_auto_out_ar_bits_echo_tl_state_size),
    .auto_out_ar_bits_echo_tl_state_source(tl2axi4_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_r_ready(tl2axi4_auto_out_r_ready),
    .auto_out_r_valid(tl2axi4_auto_out_r_valid),
    .auto_out_r_bits_id(tl2axi4_auto_out_r_bits_id),
    .auto_out_r_bits_data(tl2axi4_auto_out_r_bits_data),
    .auto_out_r_bits_resp(tl2axi4_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_tl_state_size(tl2axi4_auto_out_r_bits_echo_tl_state_size),
    .auto_out_r_bits_echo_tl_state_source(tl2axi4_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_last(tl2axi4_auto_out_r_bits_last),
    .io_covSum(tl2axi4_io_covSum),
    .metaReset(tl2axi4_metaReset)
  );
  assign widget_auto_in_a_ready = widget_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_valid = widget_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_opcode = widget_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_size = widget_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_source = widget_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_denied = widget_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_data = widget_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_corrupt = widget_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_out_a_valid = widget_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_opcode = widget_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_size = widget_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_source = widget_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_address = widget_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_bufferable = widget_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_modifiable = widget_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_readalloc = widget_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_writealloc = widget_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_privileged = widget_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_secure = widget_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_fetch = widget_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_mask = widget_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_data = widget_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_d_ready = widget_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_axi4yank_out_aw_valid = axi4yank_auto_out_aw_valid; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_aw_bits_id = axi4yank_auto_out_aw_bits_id; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_aw_bits_addr = axi4yank_auto_out_aw_bits_addr; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_aw_bits_len = axi4yank_auto_out_aw_bits_len; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_aw_bits_size = axi4yank_auto_out_aw_bits_size; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_aw_bits_burst = axi4yank_auto_out_aw_bits_burst; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_aw_bits_lock = axi4yank_auto_out_aw_bits_lock; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_aw_bits_cache = axi4yank_auto_out_aw_bits_cache; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_aw_bits_prot = axi4yank_auto_out_aw_bits_prot; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_aw_bits_qos = axi4yank_auto_out_aw_bits_qos; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_w_valid = axi4yank_auto_out_w_valid; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_w_bits_data = axi4yank_auto_out_w_bits_data; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_w_bits_strb = axi4yank_auto_out_w_bits_strb; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_w_bits_last = axi4yank_auto_out_w_bits_last; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_b_ready = axi4yank_auto_out_b_ready; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_valid = axi4yank_auto_out_ar_valid; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_bits_id = axi4yank_auto_out_ar_bits_id; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_bits_addr = axi4yank_auto_out_ar_bits_addr; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_bits_len = axi4yank_auto_out_ar_bits_len; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_bits_size = axi4yank_auto_out_ar_bits_size; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_bits_burst = axi4yank_auto_out_ar_bits_burst; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_bits_lock = axi4yank_auto_out_ar_bits_lock; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_bits_cache = axi4yank_auto_out_ar_bits_cache; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_bits_prot = axi4yank_auto_out_ar_bits_prot; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_ar_bits_qos = axi4yank_auto_out_ar_bits_qos; // @[LazyModule.scala 311:12]
  assign auto_axi4yank_out_r_ready = axi4yank_auto_out_r_ready; // @[LazyModule.scala 311:12]
  assign auto_tl_in_a_ready = widget_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_valid = widget_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_opcode = widget_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_size = widget_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_source = widget_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_denied = widget_auto_in_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_data = widget_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_tl_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign axi4yank_clock = clock;
  assign axi4yank_reset = reset;
  assign axi4yank_auto_in_aw_valid = axi4index_auto_out_aw_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_id = axi4index_auto_out_aw_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_addr = axi4index_auto_out_aw_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_len = axi4index_auto_out_aw_bits_len; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_size = axi4index_auto_out_aw_bits_size; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_burst = axi4index_auto_out_aw_bits_burst; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_lock = axi4index_auto_out_aw_bits_lock; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_cache = axi4index_auto_out_aw_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_prot = axi4index_auto_out_aw_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_qos = axi4index_auto_out_aw_bits_qos; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_echo_tl_state_size = axi4index_auto_out_aw_bits_echo_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_echo_tl_state_source = axi4index_auto_out_aw_bits_echo_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_echo_extra_id = axi4index_auto_out_aw_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_valid = axi4index_auto_out_w_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_bits_data = axi4index_auto_out_w_bits_data; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_bits_strb = axi4index_auto_out_w_bits_strb; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_bits_last = axi4index_auto_out_w_bits_last; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_b_ready = axi4index_auto_out_b_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_valid = axi4index_auto_out_ar_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_id = axi4index_auto_out_ar_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_addr = axi4index_auto_out_ar_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_len = axi4index_auto_out_ar_bits_len; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_size = axi4index_auto_out_ar_bits_size; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_burst = axi4index_auto_out_ar_bits_burst; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_lock = axi4index_auto_out_ar_bits_lock; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_cache = axi4index_auto_out_ar_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_prot = axi4index_auto_out_ar_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_qos = axi4index_auto_out_ar_bits_qos; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_echo_tl_state_size = axi4index_auto_out_ar_bits_echo_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_echo_tl_state_source = axi4index_auto_out_ar_bits_echo_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_echo_extra_id = axi4index_auto_out_ar_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_r_ready = axi4index_auto_out_r_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_aw_ready = auto_axi4yank_out_aw_ready; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_w_ready = auto_axi4yank_out_w_ready; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_b_valid = auto_axi4yank_out_b_valid; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_b_bits_id = auto_axi4yank_out_b_bits_id; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_b_bits_resp = auto_axi4yank_out_b_bits_resp; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_ar_ready = auto_axi4yank_out_ar_ready; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_r_valid = auto_axi4yank_out_r_valid; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_r_bits_id = auto_axi4yank_out_r_bits_id; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_r_bits_data = auto_axi4yank_out_r_bits_data; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_r_bits_resp = auto_axi4yank_out_r_bits_resp; // @[LazyModule.scala 311:12]
  assign axi4yank_auto_out_r_bits_last = auto_axi4yank_out_r_bits_last; // @[LazyModule.scala 311:12]
  assign axi4index_auto_in_aw_valid = tl2axi4_auto_out_aw_valid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_id = tl2axi4_auto_out_aw_bits_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_addr = tl2axi4_auto_out_aw_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_len = tl2axi4_auto_out_aw_bits_len; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_size = tl2axi4_auto_out_aw_bits_size; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_burst = tl2axi4_auto_out_aw_bits_burst; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_lock = tl2axi4_auto_out_aw_bits_lock; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_cache = tl2axi4_auto_out_aw_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_prot = tl2axi4_auto_out_aw_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_qos = tl2axi4_auto_out_aw_bits_qos; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_echo_tl_state_size = tl2axi4_auto_out_aw_bits_echo_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_aw_bits_echo_tl_state_source = tl2axi4_auto_out_aw_bits_echo_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_w_valid = tl2axi4_auto_out_w_valid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_w_bits_data = tl2axi4_auto_out_w_bits_data; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_w_bits_strb = tl2axi4_auto_out_w_bits_strb; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_w_bits_last = tl2axi4_auto_out_w_bits_last; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_b_ready = tl2axi4_auto_out_b_ready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_valid = tl2axi4_auto_out_ar_valid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_id = tl2axi4_auto_out_ar_bits_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_addr = tl2axi4_auto_out_ar_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_len = tl2axi4_auto_out_ar_bits_len; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_size = tl2axi4_auto_out_ar_bits_size; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_burst = tl2axi4_auto_out_ar_bits_burst; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_lock = tl2axi4_auto_out_ar_bits_lock; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_cache = tl2axi4_auto_out_ar_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_prot = tl2axi4_auto_out_ar_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_qos = tl2axi4_auto_out_ar_bits_qos; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_echo_tl_state_size = tl2axi4_auto_out_ar_bits_echo_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_ar_bits_echo_tl_state_source = tl2axi4_auto_out_ar_bits_echo_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4index_auto_in_r_ready = tl2axi4_auto_out_r_ready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_aw_ready = axi4yank_auto_in_aw_ready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_w_ready = axi4yank_auto_in_w_ready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_valid = axi4yank_auto_in_b_valid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_bits_id = axi4yank_auto_in_b_bits_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_bits_resp = axi4yank_auto_in_b_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_bits_echo_tl_state_size = axi4yank_auto_in_b_bits_echo_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_bits_echo_tl_state_source = axi4yank_auto_in_b_bits_echo_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_b_bits_echo_extra_id = axi4yank_auto_in_b_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_ar_ready = axi4yank_auto_in_ar_ready; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_valid = axi4yank_auto_in_r_valid; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_id = axi4yank_auto_in_r_bits_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_data = axi4yank_auto_in_r_bits_data; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_resp = axi4yank_auto_in_r_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_echo_tl_state_size = axi4yank_auto_in_r_bits_echo_tl_state_size; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_echo_tl_state_source = axi4yank_auto_in_r_bits_echo_tl_state_source; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_echo_extra_id = axi4yank_auto_in_r_bits_echo_extra_id; // @[LazyModule.scala 296:16]
  assign axi4index_auto_out_r_bits_last = axi4yank_auto_in_r_bits_last; // @[LazyModule.scala 296:16]
  assign tl2axi4_clock = clock;
  assign tl2axi4_reset = reset;
  assign tl2axi4_auto_in_a_valid = widget_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_size = widget_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_source = widget_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_address = widget_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_user_amba_prot_bufferable = widget_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_user_amba_prot_modifiable = widget_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_user_amba_prot_readalloc = widget_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_user_amba_prot_writealloc = widget_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_user_amba_prot_privileged = widget_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_user_amba_prot_secure = widget_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_user_amba_prot_fetch = widget_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_mask = widget_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_a_bits_data = widget_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_in_d_ready = widget_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_aw_ready = axi4index_auto_in_aw_ready; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_w_ready = axi4index_auto_in_w_ready; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_b_valid = axi4index_auto_in_b_valid; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_b_bits_id = axi4index_auto_in_b_bits_id; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_b_bits_resp = axi4index_auto_in_b_bits_resp; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_b_bits_echo_tl_state_size = axi4index_auto_in_b_bits_echo_tl_state_size; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_b_bits_echo_tl_state_source = axi4index_auto_in_b_bits_echo_tl_state_source; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_ar_ready = axi4index_auto_in_ar_ready; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_r_valid = axi4index_auto_in_r_valid; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_r_bits_id = axi4index_auto_in_r_bits_id; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_r_bits_data = axi4index_auto_in_r_bits_data; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_r_bits_resp = axi4index_auto_in_r_bits_resp; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_r_bits_echo_tl_state_size = axi4index_auto_in_r_bits_echo_tl_state_size; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_r_bits_echo_tl_state_source = axi4index_auto_in_r_bits_echo_tl_state_source; // @[LazyModule.scala 296:16]
  assign tl2axi4_auto_out_r_bits_last = axi4index_auto_in_r_bits_last; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_valid = auto_tl_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_opcode = auto_tl_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_size = auto_tl_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_source = auto_tl_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_address = auto_tl_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_user_amba_prot_bufferable = auto_tl_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_user_amba_prot_modifiable = auto_tl_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_user_amba_prot_readalloc = auto_tl_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_user_amba_prot_writealloc = auto_tl_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_user_amba_prot_privileged = auto_tl_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_user_amba_prot_secure = auto_tl_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_user_amba_prot_fetch = auto_tl_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_mask = auto_tl_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_bits_data = auto_tl_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_d_ready = auto_tl_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_ready = tl2axi4_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_valid = tl2axi4_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_opcode = tl2axi4_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_size = tl2axi4_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_source = tl2axi4_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_denied = tl2axi4_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_data = tl2axi4_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_corrupt = tl2axi4_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign TLInterconnectCoupler_13_covSum = 30'h0;
  assign axi4yank_sum = TLInterconnectCoupler_13_covSum + axi4yank_io_covSum;
  assign axi4index_sum = axi4yank_sum + axi4index_io_covSum;
  assign tl2axi4_sum = axi4index_sum + tl2axi4_io_covSum;
  assign io_covSum = tl2axi4_sum;
  assign tl2axi4_metaReset = metaReset;
endmodule
module MemoryBus(
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id,
  output [31:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr,
  output [7:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len,
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size,
  output [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_lock,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_cache,
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_prot,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_qos,
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid,
  output [63:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data,
  output [7:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready,
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid,
  input  [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id,
  input  [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp,
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id,
  output [31:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr,
  output [7:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len,
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size,
  output [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_lock,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_cache,
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_prot,
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_qos,
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready,
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid,
  input  [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id,
  input  [63:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data,
  input  [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp,
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last,
  input         auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock,
  input         auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset,
  output        auto_bus_xing_in_a_ready,
  input         auto_bus_xing_in_a_valid,
  input  [2:0]  auto_bus_xing_in_a_bits_opcode,
  input  [2:0]  auto_bus_xing_in_a_bits_size,
  input  [8:0]  auto_bus_xing_in_a_bits_source,
  input  [31:0] auto_bus_xing_in_a_bits_address,
  input         auto_bus_xing_in_a_bits_user_amba_prot_bufferable,
  input         auto_bus_xing_in_a_bits_user_amba_prot_modifiable,
  input         auto_bus_xing_in_a_bits_user_amba_prot_readalloc,
  input         auto_bus_xing_in_a_bits_user_amba_prot_writealloc,
  input         auto_bus_xing_in_a_bits_user_amba_prot_privileged,
  input         auto_bus_xing_in_a_bits_user_amba_prot_secure,
  input         auto_bus_xing_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_bus_xing_in_a_bits_mask,
  input  [63:0] auto_bus_xing_in_a_bits_data,
  input         auto_bus_xing_in_d_ready,
  output        auto_bus_xing_in_d_valid,
  output [2:0]  auto_bus_xing_in_d_bits_opcode,
  output [2:0]  auto_bus_xing_in_d_bits_size,
  output [8:0]  auto_bus_xing_in_d_bits_source,
  output        auto_bus_xing_in_d_bits_denied,
  output [63:0] auto_bus_xing_in_d_bits_data,
  output        auto_bus_xing_in_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_clock;
  wire  subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_reset;
  wire  subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_clock;
  wire  subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_reset;
  wire  clockGroup_auto_in_member_subsystem_mbus_0_clock;
  wire  clockGroup_auto_in_member_subsystem_mbus_0_reset;
  wire  clockGroup_auto_out_clock;
  wire  clockGroup_auto_out_reset;
  wire  fixedClockNode_auto_in_clock;
  wire  fixedClockNode_auto_in_reset;
  wire  fixedClockNode_auto_out_clock;
  wire  fixedClockNode_auto_out_reset;
  wire  subsystem_mbus_xbar_auto_in_a_ready;
  wire  subsystem_mbus_xbar_auto_in_a_valid;
  wire [2:0] subsystem_mbus_xbar_auto_in_a_bits_opcode;
  wire [2:0] subsystem_mbus_xbar_auto_in_a_bits_size;
  wire [8:0] subsystem_mbus_xbar_auto_in_a_bits_source;
  wire [31:0] subsystem_mbus_xbar_auto_in_a_bits_address;
  wire  subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_bufferable;
  wire  subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_modifiable;
  wire  subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_readalloc;
  wire  subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_writealloc;
  wire  subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_privileged;
  wire  subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_secure;
  wire  subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] subsystem_mbus_xbar_auto_in_a_bits_mask;
  wire [63:0] subsystem_mbus_xbar_auto_in_a_bits_data;
  wire  subsystem_mbus_xbar_auto_in_d_ready;
  wire  subsystem_mbus_xbar_auto_in_d_valid;
  wire [2:0] subsystem_mbus_xbar_auto_in_d_bits_opcode;
  wire [2:0] subsystem_mbus_xbar_auto_in_d_bits_size;
  wire [8:0] subsystem_mbus_xbar_auto_in_d_bits_source;
  wire  subsystem_mbus_xbar_auto_in_d_bits_denied;
  wire [63:0] subsystem_mbus_xbar_auto_in_d_bits_data;
  wire  subsystem_mbus_xbar_auto_in_d_bits_corrupt;
  wire  subsystem_mbus_xbar_auto_out_a_ready;
  wire  subsystem_mbus_xbar_auto_out_a_valid;
  wire [2:0] subsystem_mbus_xbar_auto_out_a_bits_opcode;
  wire [2:0] subsystem_mbus_xbar_auto_out_a_bits_size;
  wire [8:0] subsystem_mbus_xbar_auto_out_a_bits_source;
  wire [31:0] subsystem_mbus_xbar_auto_out_a_bits_address;
  wire  subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_bufferable;
  wire  subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_modifiable;
  wire  subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_readalloc;
  wire  subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_writealloc;
  wire  subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_privileged;
  wire  subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_secure;
  wire  subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] subsystem_mbus_xbar_auto_out_a_bits_mask;
  wire [63:0] subsystem_mbus_xbar_auto_out_a_bits_data;
  wire  subsystem_mbus_xbar_auto_out_d_ready;
  wire  subsystem_mbus_xbar_auto_out_d_valid;
  wire [2:0] subsystem_mbus_xbar_auto_out_d_bits_opcode;
  wire [2:0] subsystem_mbus_xbar_auto_out_d_bits_size;
  wire [8:0] subsystem_mbus_xbar_auto_out_d_bits_source;
  wire  subsystem_mbus_xbar_auto_out_d_bits_denied;
  wire [63:0] subsystem_mbus_xbar_auto_out_d_bits_data;
  wire  subsystem_mbus_xbar_auto_out_d_bits_corrupt;
  wire  fixer_auto_in_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [8:0] fixer_auto_in_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_in_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_in_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [8:0] fixer_auto_in_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [8:0] fixer_auto_out_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_out_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_out_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [8:0] fixer_auto_out_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire [29:0] fixer_io_covSum; // @[FIFOFixer.scala 144:27]
  wire  picker_auto_in_a_ready; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_a_valid; // @[ProbePicker.scala 65:28]
  wire [2:0] picker_auto_in_a_bits_opcode; // @[ProbePicker.scala 65:28]
  wire [2:0] picker_auto_in_a_bits_size; // @[ProbePicker.scala 65:28]
  wire [8:0] picker_auto_in_a_bits_source; // @[ProbePicker.scala 65:28]
  wire [31:0] picker_auto_in_a_bits_address; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_a_bits_user_amba_prot_bufferable; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_a_bits_user_amba_prot_modifiable; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_a_bits_user_amba_prot_readalloc; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_a_bits_user_amba_prot_writealloc; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_a_bits_user_amba_prot_privileged; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_a_bits_user_amba_prot_secure; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_a_bits_user_amba_prot_fetch; // @[ProbePicker.scala 65:28]
  wire [7:0] picker_auto_in_a_bits_mask; // @[ProbePicker.scala 65:28]
  wire [63:0] picker_auto_in_a_bits_data; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_d_ready; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_d_valid; // @[ProbePicker.scala 65:28]
  wire [2:0] picker_auto_in_d_bits_opcode; // @[ProbePicker.scala 65:28]
  wire [2:0] picker_auto_in_d_bits_size; // @[ProbePicker.scala 65:28]
  wire [8:0] picker_auto_in_d_bits_source; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_d_bits_denied; // @[ProbePicker.scala 65:28]
  wire [63:0] picker_auto_in_d_bits_data; // @[ProbePicker.scala 65:28]
  wire  picker_auto_in_d_bits_corrupt; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_a_ready; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_a_valid; // @[ProbePicker.scala 65:28]
  wire [2:0] picker_auto_out_a_bits_opcode; // @[ProbePicker.scala 65:28]
  wire [2:0] picker_auto_out_a_bits_size; // @[ProbePicker.scala 65:28]
  wire [8:0] picker_auto_out_a_bits_source; // @[ProbePicker.scala 65:28]
  wire [31:0] picker_auto_out_a_bits_address; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_a_bits_user_amba_prot_bufferable; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_a_bits_user_amba_prot_modifiable; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_a_bits_user_amba_prot_readalloc; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_a_bits_user_amba_prot_writealloc; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_a_bits_user_amba_prot_privileged; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_a_bits_user_amba_prot_secure; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_a_bits_user_amba_prot_fetch; // @[ProbePicker.scala 65:28]
  wire [7:0] picker_auto_out_a_bits_mask; // @[ProbePicker.scala 65:28]
  wire [63:0] picker_auto_out_a_bits_data; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_d_ready; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_d_valid; // @[ProbePicker.scala 65:28]
  wire [2:0] picker_auto_out_d_bits_opcode; // @[ProbePicker.scala 65:28]
  wire [2:0] picker_auto_out_d_bits_size; // @[ProbePicker.scala 65:28]
  wire [8:0] picker_auto_out_d_bits_source; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_d_bits_denied; // @[ProbePicker.scala 65:28]
  wire [63:0] picker_auto_out_d_bits_data; // @[ProbePicker.scala 65:28]
  wire  picker_auto_out_d_bits_corrupt; // @[ProbePicker.scala 65:28]
  wire [29:0] picker_io_covSum; // @[ProbePicker.scala 65:28]
  wire  buffer_auto_in_a_ready;
  wire  buffer_auto_in_a_valid;
  wire [2:0] buffer_auto_in_a_bits_opcode;
  wire [2:0] buffer_auto_in_a_bits_size;
  wire [8:0] buffer_auto_in_a_bits_source;
  wire [31:0] buffer_auto_in_a_bits_address;
  wire  buffer_auto_in_a_bits_user_amba_prot_bufferable;
  wire  buffer_auto_in_a_bits_user_amba_prot_modifiable;
  wire  buffer_auto_in_a_bits_user_amba_prot_readalloc;
  wire  buffer_auto_in_a_bits_user_amba_prot_writealloc;
  wire  buffer_auto_in_a_bits_user_amba_prot_privileged;
  wire  buffer_auto_in_a_bits_user_amba_prot_secure;
  wire  buffer_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] buffer_auto_in_a_bits_mask;
  wire [63:0] buffer_auto_in_a_bits_data;
  wire  buffer_auto_in_d_ready;
  wire  buffer_auto_in_d_valid;
  wire [2:0] buffer_auto_in_d_bits_opcode;
  wire [2:0] buffer_auto_in_d_bits_size;
  wire [8:0] buffer_auto_in_d_bits_source;
  wire  buffer_auto_in_d_bits_denied;
  wire [63:0] buffer_auto_in_d_bits_data;
  wire  buffer_auto_in_d_bits_corrupt;
  wire  buffer_auto_out_a_ready;
  wire  buffer_auto_out_a_valid;
  wire [2:0] buffer_auto_out_a_bits_opcode;
  wire [2:0] buffer_auto_out_a_bits_size;
  wire [8:0] buffer_auto_out_a_bits_source;
  wire [31:0] buffer_auto_out_a_bits_address;
  wire  buffer_auto_out_a_bits_user_amba_prot_bufferable;
  wire  buffer_auto_out_a_bits_user_amba_prot_modifiable;
  wire  buffer_auto_out_a_bits_user_amba_prot_readalloc;
  wire  buffer_auto_out_a_bits_user_amba_prot_writealloc;
  wire  buffer_auto_out_a_bits_user_amba_prot_privileged;
  wire  buffer_auto_out_a_bits_user_amba_prot_secure;
  wire  buffer_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] buffer_auto_out_a_bits_mask;
  wire [63:0] buffer_auto_out_a_bits_data;
  wire  buffer_auto_out_d_ready;
  wire  buffer_auto_out_d_valid;
  wire [2:0] buffer_auto_out_d_bits_opcode;
  wire [2:0] buffer_auto_out_d_bits_size;
  wire [8:0] buffer_auto_out_d_bits_source;
  wire  buffer_auto_out_d_bits_denied;
  wire [63:0] buffer_auto_out_d_bits_data;
  wire  buffer_auto_out_d_bits_corrupt;
  wire  coupler_to_memory_controller_port_named_axi4_clock; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_reset; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_valid; // @[LazyModule.scala 432:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_id; // @[LazyModule.scala 432:27]
  wire [31:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_addr; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_len; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_size; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_burst; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_lock; // @[LazyModule.scala 432:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_cache; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_prot; // @[LazyModule.scala 432:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_qos; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_valid; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_data; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_strb; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_last; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_valid; // @[LazyModule.scala 432:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_id; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_resp; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_valid; // @[LazyModule.scala 432:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_id; // @[LazyModule.scala 432:27]
  wire [31:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_addr; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_len; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_size; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_burst; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_lock; // @[LazyModule.scala 432:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_cache; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_prot; // @[LazyModule.scala 432:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_qos; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_valid; // @[LazyModule.scala 432:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_id; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_data; // @[LazyModule.scala 432:27]
  wire [1:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_resp; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_last; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_size; // @[LazyModule.scala 432:27]
  wire [8:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_source; // @[LazyModule.scala 432:27]
  wire [31:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_address; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_secure; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 432:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_mask; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_ready; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size; // @[LazyModule.scala 432:27]
  wire [8:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied; // @[LazyModule.scala 432:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_data; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt; // @[LazyModule.scala 432:27]
  wire [29:0] coupler_to_memory_controller_port_named_axi4_io_covSum; // @[LazyModule.scala 432:27]
  wire  coupler_to_memory_controller_port_named_axi4_metaReset; // @[LazyModule.scala 432:27]
  wire [29:0] MemoryBus_covSum;
  wire [29:0] fixer_sum;
  wire [29:0] picker_sum;
  wire [29:0] coupler_to_memory_controller_port_named_axi4_sum;
  TLFIFOFixer_4 fixer ( // @[FIFOFixer.scala 144:27]
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(fixer_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(fixer_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(fixer_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(fixer_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(fixer_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(fixer_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(fixer_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_auto_in_a_bits_data),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(fixer_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(fixer_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(fixer_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(fixer_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(fixer_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(fixer_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(fixer_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_auto_out_a_bits_data),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt),
    .io_covSum(fixer_io_covSum)
  );
  ProbePicker picker ( // @[ProbePicker.scala 65:28]
    .auto_in_a_ready(picker_auto_in_a_ready),
    .auto_in_a_valid(picker_auto_in_a_valid),
    .auto_in_a_bits_opcode(picker_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(picker_auto_in_a_bits_size),
    .auto_in_a_bits_source(picker_auto_in_a_bits_source),
    .auto_in_a_bits_address(picker_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(picker_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(picker_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(picker_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(picker_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(picker_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(picker_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(picker_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(picker_auto_in_a_bits_mask),
    .auto_in_a_bits_data(picker_auto_in_a_bits_data),
    .auto_in_d_ready(picker_auto_in_d_ready),
    .auto_in_d_valid(picker_auto_in_d_valid),
    .auto_in_d_bits_opcode(picker_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(picker_auto_in_d_bits_size),
    .auto_in_d_bits_source(picker_auto_in_d_bits_source),
    .auto_in_d_bits_denied(picker_auto_in_d_bits_denied),
    .auto_in_d_bits_data(picker_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(picker_auto_in_d_bits_corrupt),
    .auto_out_a_ready(picker_auto_out_a_ready),
    .auto_out_a_valid(picker_auto_out_a_valid),
    .auto_out_a_bits_opcode(picker_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(picker_auto_out_a_bits_size),
    .auto_out_a_bits_source(picker_auto_out_a_bits_source),
    .auto_out_a_bits_address(picker_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(picker_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(picker_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(picker_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(picker_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(picker_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(picker_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(picker_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(picker_auto_out_a_bits_mask),
    .auto_out_a_bits_data(picker_auto_out_a_bits_data),
    .auto_out_d_ready(picker_auto_out_d_ready),
    .auto_out_d_valid(picker_auto_out_d_valid),
    .auto_out_d_bits_opcode(picker_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(picker_auto_out_d_bits_size),
    .auto_out_d_bits_source(picker_auto_out_d_bits_source),
    .auto_out_d_bits_denied(picker_auto_out_d_bits_denied),
    .auto_out_d_bits_data(picker_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(picker_auto_out_d_bits_corrupt),
    .io_covSum(picker_io_covSum)
  );
  TLInterconnectCoupler_13 coupler_to_memory_controller_port_named_axi4 ( // @[LazyModule.scala 432:27]
    .clock(coupler_to_memory_controller_port_named_axi4_clock),
    .reset(coupler_to_memory_controller_port_named_axi4_reset),
    .auto_axi4yank_out_aw_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_ready),
    .auto_axi4yank_out_aw_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_valid),
    .auto_axi4yank_out_aw_bits_id(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_id),
    .auto_axi4yank_out_aw_bits_addr(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_addr),
    .auto_axi4yank_out_aw_bits_len(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_len),
    .auto_axi4yank_out_aw_bits_size(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_size),
    .auto_axi4yank_out_aw_bits_burst(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_burst),
    .auto_axi4yank_out_aw_bits_lock(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_lock),
    .auto_axi4yank_out_aw_bits_cache(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_cache),
    .auto_axi4yank_out_aw_bits_prot(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_prot),
    .auto_axi4yank_out_aw_bits_qos(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_qos),
    .auto_axi4yank_out_w_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_ready),
    .auto_axi4yank_out_w_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_valid),
    .auto_axi4yank_out_w_bits_data(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_data),
    .auto_axi4yank_out_w_bits_strb(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_strb),
    .auto_axi4yank_out_w_bits_last(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_last),
    .auto_axi4yank_out_b_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_ready),
    .auto_axi4yank_out_b_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_valid),
    .auto_axi4yank_out_b_bits_id(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_id),
    .auto_axi4yank_out_b_bits_resp(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_resp),
    .auto_axi4yank_out_ar_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_ready),
    .auto_axi4yank_out_ar_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_valid),
    .auto_axi4yank_out_ar_bits_id(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_id),
    .auto_axi4yank_out_ar_bits_addr(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_addr),
    .auto_axi4yank_out_ar_bits_len(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_len),
    .auto_axi4yank_out_ar_bits_size(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_size),
    .auto_axi4yank_out_ar_bits_burst(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_burst),
    .auto_axi4yank_out_ar_bits_lock(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_lock),
    .auto_axi4yank_out_ar_bits_cache(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_cache),
    .auto_axi4yank_out_ar_bits_prot(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_prot),
    .auto_axi4yank_out_ar_bits_qos(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_qos),
    .auto_axi4yank_out_r_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_ready),
    .auto_axi4yank_out_r_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_valid),
    .auto_axi4yank_out_r_bits_id(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_id),
    .auto_axi4yank_out_r_bits_data(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_data),
    .auto_axi4yank_out_r_bits_resp(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_resp),
    .auto_axi4yank_out_r_bits_last(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_last),
    .auto_tl_in_a_ready(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready),
    .auto_tl_in_a_valid(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_valid),
    .auto_tl_in_a_bits_opcode(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_opcode),
    .auto_tl_in_a_bits_size(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_size),
    .auto_tl_in_a_bits_source(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_source),
    .auto_tl_in_a_bits_address(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_address),
    .auto_tl_in_a_bits_user_amba_prot_bufferable(
      coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_bufferable),
    .auto_tl_in_a_bits_user_amba_prot_modifiable(
      coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_modifiable),
    .auto_tl_in_a_bits_user_amba_prot_readalloc(
      coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_readalloc),
    .auto_tl_in_a_bits_user_amba_prot_writealloc(
      coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_writealloc),
    .auto_tl_in_a_bits_user_amba_prot_privileged(
      coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_privileged),
    .auto_tl_in_a_bits_user_amba_prot_secure(
      coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_secure),
    .auto_tl_in_a_bits_user_amba_prot_fetch(
      coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_fetch),
    .auto_tl_in_a_bits_mask(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_mask),
    .auto_tl_in_a_bits_data(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_data),
    .auto_tl_in_d_ready(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_ready),
    .auto_tl_in_d_valid(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_opcode(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode),
    .auto_tl_in_d_bits_size(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_denied(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied),
    .auto_tl_in_d_bits_data(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_data),
    .auto_tl_in_d_bits_corrupt(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt),
    .io_covSum(coupler_to_memory_controller_port_named_axi4_io_covSum),
    .metaReset(coupler_to_memory_controller_port_named_axi4_metaReset)
  );
  assign subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_clock =
    subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_reset =
    subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_clock = clockGroup_auto_in_member_subsystem_mbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_reset = clockGroup_auto_in_member_subsystem_mbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fixedClockNode_auto_out_clock = fixedClockNode_auto_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fixedClockNode_auto_out_reset = fixedClockNode_auto_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_in_a_ready = subsystem_mbus_xbar_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_mbus_xbar_auto_in_d_valid = subsystem_mbus_xbar_auto_out_d_valid; // @[ReadyValidCancel.scala 21:38]
  assign subsystem_mbus_xbar_auto_in_d_bits_opcode = subsystem_mbus_xbar_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_mbus_xbar_auto_in_d_bits_size = subsystem_mbus_xbar_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_mbus_xbar_auto_in_d_bits_source = subsystem_mbus_xbar_auto_out_d_bits_source; // @[Xbar.scala 228:69]
  assign subsystem_mbus_xbar_auto_in_d_bits_denied = subsystem_mbus_xbar_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_mbus_xbar_auto_in_d_bits_data = subsystem_mbus_xbar_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_mbus_xbar_auto_in_d_bits_corrupt = subsystem_mbus_xbar_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_mbus_xbar_auto_out_a_valid = subsystem_mbus_xbar_auto_in_a_valid; // @[ReadyValidCancel.scala 21:38]
  assign subsystem_mbus_xbar_auto_out_a_bits_opcode = subsystem_mbus_xbar_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_size = subsystem_mbus_xbar_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_source = subsystem_mbus_xbar_auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign subsystem_mbus_xbar_auto_out_a_bits_address = subsystem_mbus_xbar_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_bufferable =
    subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_modifiable =
    subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_readalloc =
    subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_writealloc =
    subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_privileged =
    subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_secure =
    subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_fetch =
    subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_mask = subsystem_mbus_xbar_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_a_bits_data = subsystem_mbus_xbar_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_mbus_xbar_auto_out_d_ready = subsystem_mbus_xbar_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_ready = buffer_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_valid = buffer_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_opcode = buffer_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_size = buffer_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_source = buffer_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_denied = buffer_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_data = buffer_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_corrupt = buffer_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_a_valid = buffer_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_opcode = buffer_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_size = buffer_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_source = buffer_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_address = buffer_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_bufferable = buffer_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_modifiable = buffer_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_readalloc = buffer_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_writealloc = buffer_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_privileged = buffer_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_secure = buffer_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_fetch = buffer_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_mask = buffer_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_data = buffer_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_d_ready = buffer_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_id; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_addr; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_len; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_burst; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_lock =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_lock; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_cache =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_cache; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_prot =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_prot; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_qos =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_qos; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_data; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_strb; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_last; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_ready; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_id; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_addr; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_len; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_burst; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_lock =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_lock; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_cache =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_cache; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_prot =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_prot; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_qos =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_qos; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_ready; // @[LazyModule.scala 311:12]
  assign auto_bus_xing_in_a_ready = buffer_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_valid = buffer_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_size = buffer_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_source = buffer_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_denied = buffer_auto_in_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_data = buffer_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_bus_xing_in_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_clock =
    auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock; // @[LazyModule.scala 309:16]
  assign subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_reset =
    auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset; // @[LazyModule.scala 309:16]
  assign clockGroup_auto_in_member_subsystem_mbus_0_clock =
    subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_clock; // @[LazyModule.scala 298:16]
  assign clockGroup_auto_in_member_subsystem_mbus_0_reset =
    subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_reset; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[LazyModule.scala 298:16]
  assign subsystem_mbus_xbar_auto_in_a_valid = fixer_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_size = fixer_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_source = fixer_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_address = fixer_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_bufferable = fixer_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_modifiable = fixer_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_readalloc = fixer_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_writealloc = fixer_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_privileged = fixer_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_secure = fixer_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_user_amba_prot_fetch = fixer_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_a_bits_data = fixer_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_in_d_ready = fixer_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_xbar_auto_out_a_ready = picker_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_mbus_xbar_auto_out_d_valid = picker_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_mbus_xbar_auto_out_d_bits_opcode = picker_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_mbus_xbar_auto_out_d_bits_size = picker_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_mbus_xbar_auto_out_d_bits_source = picker_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_mbus_xbar_auto_out_d_bits_denied = picker_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign subsystem_mbus_xbar_auto_out_d_bits_data = picker_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_mbus_xbar_auto_out_d_bits_corrupt = picker_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign fixer_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_bufferable = buffer_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_modifiable = buffer_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_readalloc = buffer_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_writealloc = buffer_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_privileged = buffer_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_secure = buffer_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_fetch = buffer_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_a_ready = subsystem_mbus_xbar_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_valid = subsystem_mbus_xbar_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_opcode = subsystem_mbus_xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_size = subsystem_mbus_xbar_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_source = subsystem_mbus_xbar_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_denied = subsystem_mbus_xbar_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_data = subsystem_mbus_xbar_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_corrupt = subsystem_mbus_xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign picker_auto_in_a_valid = subsystem_mbus_xbar_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_opcode = subsystem_mbus_xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_size = subsystem_mbus_xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_source = subsystem_mbus_xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_address = subsystem_mbus_xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_user_amba_prot_bufferable = subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_bufferable
    ; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_user_amba_prot_modifiable = subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_modifiable
    ; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_user_amba_prot_readalloc = subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_user_amba_prot_writealloc = subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_writealloc
    ; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_user_amba_prot_privileged = subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_privileged
    ; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_user_amba_prot_secure = subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_user_amba_prot_fetch = subsystem_mbus_xbar_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_mask = subsystem_mbus_xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign picker_auto_in_a_bits_data = subsystem_mbus_xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign picker_auto_in_d_ready = subsystem_mbus_xbar_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign picker_auto_out_a_ready = coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready; // @[LazyModule.scala 298:16]
  assign picker_auto_out_d_valid = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid; // @[LazyModule.scala 298:16]
  assign picker_auto_out_d_bits_opcode = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign picker_auto_out_d_bits_size = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign picker_auto_out_d_bits_source = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign picker_auto_out_d_bits_denied = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign picker_auto_out_d_bits_data = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign picker_auto_out_d_bits_corrupt = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_valid = auto_bus_xing_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_opcode = auto_bus_xing_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_size = auto_bus_xing_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_source = auto_bus_xing_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_address = auto_bus_xing_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_user_amba_prot_bufferable = auto_bus_xing_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_user_amba_prot_modifiable = auto_bus_xing_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_user_amba_prot_readalloc = auto_bus_xing_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_user_amba_prot_writealloc = auto_bus_xing_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_user_amba_prot_privileged = auto_bus_xing_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_user_amba_prot_secure = auto_bus_xing_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_user_amba_prot_fetch = auto_bus_xing_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_mask = auto_bus_xing_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_data = auto_bus_xing_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_d_ready = auto_bus_xing_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_ready = fixer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_valid = fixer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_size = fixer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_source = fixer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_denied = fixer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_data = fixer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign coupler_to_memory_controller_port_named_axi4_clock = fixedClockNode_auto_out_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_memory_controller_port_named_axi4_reset = fixedClockNode_auto_out_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_ready =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_ready =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_valid =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_id =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_resp =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_ready =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_valid =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_id =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_data =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_resp =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_last =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last; // @[LazyModule.scala 311:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_valid = picker_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_opcode = picker_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_size = picker_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_source = picker_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_address = picker_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_bufferable =
    picker_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_modifiable =
    picker_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_readalloc =
    picker_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_writealloc =
    picker_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_privileged =
    picker_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_secure =
    picker_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_user_amba_prot_fetch =
    picker_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_mask = picker_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_data = picker_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_ready = picker_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign MemoryBus_covSum = 30'h0;
  assign fixer_sum = MemoryBus_covSum + fixer_io_covSum;
  assign picker_sum = fixer_sum + picker_io_covSum;
  assign coupler_to_memory_controller_port_named_axi4_sum = picker_sum +
    coupler_to_memory_controller_port_named_axi4_io_covSum;
  assign io_covSum = coupler_to_memory_controller_port_named_axi4_sum;
  assign coupler_to_memory_controller_port_named_axi4_metaReset = metaReset;
endmodule
module BroadcastFilter(
  output        io_request_ready,
  input         io_request_valid,
  input         io_response_ready,
  output        io_response_valid,
  output [29:0] io_covSum
);
  wire [29:0] BroadcastFilter_covSum;
  assign io_request_ready = io_response_ready; // @[Broadcast.scala 362:20]
  assign io_response_valid = io_request_valid; // @[Broadcast.scala 363:21]
  assign BroadcastFilter_covSum = 30'h0;
  assign io_covSum = BroadcastFilter_covSum;
endmodule
module Queue_20(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram_mask [0:7]; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_mask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:7]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] value; // @[Counter.scala 62:40]
  reg [2:0] value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 78:24]
  wire [2:0] _value_T_3 = value_1 + 3'h1; // @[Counter.scala 78:24]
  wire [29:0] Queue_20_covSum;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_20_covSum = 30'h0;
  assign io_covSum = Queue_20_covSum;
  always @(posedge clock) begin
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= _value_T_1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= _value_T_3;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_mask[initvar] = _RAND_0[7:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBroadcastTracker(
  input         clock,
  input         reset,
  input         io_in_a_first,
  output        io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input         io_in_a_bits_user_amba_prot_bufferable,
  input         io_in_a_bits_user_amba_prot_modifiable,
  input         io_in_a_bits_user_amba_prot_readalloc,
  input         io_in_a_bits_user_amba_prot_writealloc,
  input         io_in_a_bits_user_amba_prot_privileged,
  input         io_in_a_bits_user_amba_prot_secure,
  input         io_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  io_in_a_bits_mask,
  input  [63:0] io_in_a_bits_data,
  input         io_out_a_ready,
  output        io_out_a_valid,
  output [2:0]  io_out_a_bits_opcode,
  output [2:0]  io_out_a_bits_size,
  output [8:0]  io_out_a_bits_source,
  output [31:0] io_out_a_bits_address,
  output        io_out_a_bits_user_amba_prot_bufferable,
  output        io_out_a_bits_user_amba_prot_modifiable,
  output        io_out_a_bits_user_amba_prot_readalloc,
  output        io_out_a_bits_user_amba_prot_writealloc,
  output        io_out_a_bits_user_amba_prot_privileged,
  output        io_out_a_bits_user_amba_prot_secure,
  output        io_out_a_bits_user_amba_prot_fetch,
  output [7:0]  io_out_a_bits_mask,
  output [63:0] io_out_a_bits_data,
  input         io_probedack,
  input         io_d_last,
  output [6:0]  io_source,
  output [25:0] io_line,
  output        io_idle,
  output        io_need_d,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  o_data_clock; // @[Decoupled.scala 361:21]
  wire  o_data_reset; // @[Decoupled.scala 361:21]
  wire  o_data_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  o_data_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [7:0] o_data_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] o_data_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  o_data_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  o_data_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [7:0] o_data_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] o_data_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [29:0] o_data_io_covSum; // @[Decoupled.scala 361:21]
  reg  got_e; // @[Broadcast.scala 423:24]
  reg  sent_d; // @[Broadcast.scala 424:24]
  reg [2:0] opcode; // @[Broadcast.scala 426:20]
  reg [2:0] size; // @[Broadcast.scala 428:20]
  reg [6:0] source; // @[Broadcast.scala 429:20]
  reg  user_amba_prot_bufferable; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_modifiable; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_readalloc; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_writealloc; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_privileged; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_secure; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_fetch; // @[Broadcast.scala 430:20]
  reg [31:0] address; // @[Broadcast.scala 432:24]
  wire  idle = got_e & sent_d; // @[Broadcast.scala 435:23]
  wire  _T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = _T & io_in_a_first; // @[Broadcast.scala 437:24]
  wire  _T_3 = ~reset; // @[Broadcast.scala 438:12]
  wire  _GEN_0 = _T & io_in_a_first ? 1'h0 : sent_d; // @[Broadcast.scala 437:42 439:13 424:24]
  wire  _GEN_2 = _T & io_in_a_first ? io_in_a_bits_opcode != 3'h6 & io_in_a_bits_opcode != 3'h7 : got_e; // @[Broadcast.scala 437:42 441:13 423:24]
  wire  _GEN_18 = io_d_last | _GEN_0; // @[Broadcast.scala 458:20 460:12]
  wire  _io_in_a_ready_T_1 = idle | ~io_in_a_first; // @[Broadcast.scala 485:26]
  wire  i_data_ready = o_data_io_enq_ready; // @[Broadcast.scala 482:20 Decoupled.scala 365:17]
  wire  acquire = opcode == 3'h6 | opcode == 3'h7; // @[Broadcast.scala 491:52]
  wire [1:0] _io_out_a_bits_source_T = acquire ? 2'h3 : 2'h0; // @[Broadcast.scala 500:35]
  wire [29:0] TLBroadcastTracker_covSum;
  wire [29:0] o_data_sum;
  Queue_20 o_data ( // @[Decoupled.scala 361:21]
    .clock(o_data_clock),
    .reset(o_data_reset),
    .io_enq_ready(o_data_io_enq_ready),
    .io_enq_valid(o_data_io_enq_valid),
    .io_enq_bits_mask(o_data_io_enq_bits_mask),
    .io_enq_bits_data(o_data_io_enq_bits_data),
    .io_deq_ready(o_data_io_deq_ready),
    .io_deq_valid(o_data_io_deq_valid),
    .io_deq_bits_mask(o_data_io_deq_bits_mask),
    .io_deq_bits_data(o_data_io_deq_bits_data),
    .io_covSum(o_data_io_covSum)
  );
  assign io_in_a_ready = (idle | ~io_in_a_first) & i_data_ready; // @[Broadcast.scala 485:45]
  assign io_out_a_valid = o_data_io_deq_valid; // @[Broadcast.scala 496:34]
  assign io_out_a_bits_opcode = acquire ? 3'h4 : opcode; // @[Broadcast.scala 497:31]
  assign io_out_a_bits_size = size; // @[Broadcast.scala 499:25]
  assign io_out_a_bits_source = {_io_out_a_bits_source_T,source}; // @[Cat.scala 31:58]
  assign io_out_a_bits_address = address; // @[Broadcast.scala 501:25]
  assign io_out_a_bits_user_amba_prot_bufferable = user_amba_prot_bufferable; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_modifiable = user_amba_prot_modifiable; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_readalloc = user_amba_prot_readalloc; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_writealloc = user_amba_prot_writealloc; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_privileged = user_amba_prot_privileged; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_secure = user_amba_prot_secure; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_fetch = user_amba_prot_fetch; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_mask = o_data_io_deq_bits_mask; // @[Broadcast.scala 502:25]
  assign io_out_a_bits_data = o_data_io_deq_bits_data; // @[Broadcast.scala 503:25]
  assign io_source = source; // @[Broadcast.scala 478:13]
  assign io_line = address[31:6]; // @[Broadcast.scala 479:22]
  assign io_idle = got_e & sent_d; // @[Broadcast.scala 435:23]
  assign io_need_d = ~sent_d; // @[Broadcast.scala 477:16]
  assign o_data_clock = clock;
  assign o_data_reset = reset;
  assign o_data_io_enq_valid = _io_in_a_ready_T_1 & io_in_a_valid; // @[Broadcast.scala 486:44]
  assign o_data_io_enq_bits_mask = io_in_a_bits_mask; // @[Broadcast.scala 482:20 487:20]
  assign o_data_io_enq_bits_data = io_in_a_bits_data; // @[Broadcast.scala 482:20 488:20]
  assign o_data_io_deq_ready = io_out_a_ready; // @[Broadcast.scala 495:34]
  assign TLBroadcastTracker_covSum = 30'h0;
  assign o_data_sum = TLBroadcastTracker_covSum + o_data_io_covSum;
  assign io_covSum = o_data_sum;
  always @(posedge clock) begin
    got_e <= reset | _GEN_2; // @[Broadcast.scala 423:{24,24}]
    sent_d <= reset | _GEN_18; // @[Broadcast.scala 424:{24,24}]
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      opcode <= io_in_a_bits_opcode; // @[Broadcast.scala 442:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      size <= io_in_a_bits_size; // @[Broadcast.scala 444:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      source <= io_in_a_bits_source; // @[Broadcast.scala 445:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_bufferable <= io_in_a_bits_user_amba_prot_bufferable; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_modifiable <= io_in_a_bits_user_amba_prot_modifiable; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_readalloc <= io_in_a_bits_user_amba_prot_readalloc; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_writealloc <= io_in_a_bits_user_amba_prot_writealloc; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_privileged <= io_in_a_bits_user_amba_prot_privileged; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_secure <= io_in_a_bits_user_amba_prot_secure; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_fetch <= io_in_a_bits_user_amba_prot_fetch; // @[BundleMap.scala 247:19]
    end
    if (reset) begin // @[Broadcast.scala 432:24]
      address <= 32'h0; // @[Broadcast.scala 432:24]
    end else if (_T & io_in_a_first) begin
      address <= io_in_a_bits_address;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~idle & (_T_1 & ~reset)) begin
          $fatal; // @[Broadcast.scala 438:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset & ~idle) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:438 assert (idle)\n"); // @[Broadcast.scala 438:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~sent_d) & (io_d_last & _T_3)) begin
          $fatal; // @[Broadcast.scala 459:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_d_last & _T_3 & ~(~sent_d)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:459 assert (!sent_d)\n"); // @[Broadcast.scala 459:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h0 & (io_probedack & _T_3)) begin
          $fatal; // @[Broadcast.scala 468:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_probedack & _T_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:468 assert (count > 0.U)\n"); // @[Broadcast.scala 468:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  got_e = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sent_d = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  opcode = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  user_amba_prot_bufferable = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  user_amba_prot_modifiable = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  user_amba_prot_readalloc = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  user_amba_prot_writealloc = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  user_amba_prot_privileged = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  user_amba_prot_secure = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  user_amba_prot_fetch = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  address = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBroadcastTracker_1(
  input         clock,
  input         reset,
  input         io_in_a_first,
  output        io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input         io_in_a_bits_user_amba_prot_bufferable,
  input         io_in_a_bits_user_amba_prot_modifiable,
  input         io_in_a_bits_user_amba_prot_readalloc,
  input         io_in_a_bits_user_amba_prot_writealloc,
  input         io_in_a_bits_user_amba_prot_privileged,
  input         io_in_a_bits_user_amba_prot_secure,
  input         io_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  io_in_a_bits_mask,
  input  [63:0] io_in_a_bits_data,
  input         io_out_a_ready,
  output        io_out_a_valid,
  output [2:0]  io_out_a_bits_opcode,
  output [2:0]  io_out_a_bits_size,
  output [8:0]  io_out_a_bits_source,
  output [31:0] io_out_a_bits_address,
  output        io_out_a_bits_user_amba_prot_bufferable,
  output        io_out_a_bits_user_amba_prot_modifiable,
  output        io_out_a_bits_user_amba_prot_readalloc,
  output        io_out_a_bits_user_amba_prot_writealloc,
  output        io_out_a_bits_user_amba_prot_privileged,
  output        io_out_a_bits_user_amba_prot_secure,
  output        io_out_a_bits_user_amba_prot_fetch,
  output [7:0]  io_out_a_bits_mask,
  output [63:0] io_out_a_bits_data,
  input         io_probedack,
  input         io_d_last,
  output [6:0]  io_source,
  output [25:0] io_line,
  output        io_idle,
  output        io_need_d,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  o_data_clock; // @[Decoupled.scala 361:21]
  wire  o_data_reset; // @[Decoupled.scala 361:21]
  wire  o_data_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  o_data_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [7:0] o_data_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] o_data_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  o_data_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  o_data_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [7:0] o_data_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] o_data_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [29:0] o_data_io_covSum; // @[Decoupled.scala 361:21]
  reg  got_e; // @[Broadcast.scala 423:24]
  reg  sent_d; // @[Broadcast.scala 424:24]
  reg [2:0] opcode; // @[Broadcast.scala 426:20]
  reg [2:0] size; // @[Broadcast.scala 428:20]
  reg [6:0] source; // @[Broadcast.scala 429:20]
  reg  user_amba_prot_bufferable; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_modifiable; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_readalloc; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_writealloc; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_privileged; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_secure; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_fetch; // @[Broadcast.scala 430:20]
  reg [31:0] address; // @[Broadcast.scala 432:24]
  wire  idle = got_e & sent_d; // @[Broadcast.scala 435:23]
  wire  _T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = _T & io_in_a_first; // @[Broadcast.scala 437:24]
  wire  _T_3 = ~reset; // @[Broadcast.scala 438:12]
  wire  _GEN_0 = _T & io_in_a_first ? 1'h0 : sent_d; // @[Broadcast.scala 437:42 439:13 424:24]
  wire  _GEN_2 = _T & io_in_a_first ? io_in_a_bits_opcode != 3'h6 & io_in_a_bits_opcode != 3'h7 : got_e; // @[Broadcast.scala 437:42 441:13 423:24]
  wire  _GEN_18 = io_d_last | _GEN_0; // @[Broadcast.scala 458:20 460:12]
  wire  _io_in_a_ready_T_1 = idle | ~io_in_a_first; // @[Broadcast.scala 485:26]
  wire  i_data_ready = o_data_io_enq_ready; // @[Broadcast.scala 482:20 Decoupled.scala 365:17]
  wire  acquire = opcode == 3'h6 | opcode == 3'h7; // @[Broadcast.scala 491:52]
  wire [1:0] _io_out_a_bits_source_T = acquire ? 2'h3 : 2'h0; // @[Broadcast.scala 500:35]
  wire [29:0] TLBroadcastTracker_1_covSum;
  wire [29:0] o_data_sum;
  Queue_20 o_data ( // @[Decoupled.scala 361:21]
    .clock(o_data_clock),
    .reset(o_data_reset),
    .io_enq_ready(o_data_io_enq_ready),
    .io_enq_valid(o_data_io_enq_valid),
    .io_enq_bits_mask(o_data_io_enq_bits_mask),
    .io_enq_bits_data(o_data_io_enq_bits_data),
    .io_deq_ready(o_data_io_deq_ready),
    .io_deq_valid(o_data_io_deq_valid),
    .io_deq_bits_mask(o_data_io_deq_bits_mask),
    .io_deq_bits_data(o_data_io_deq_bits_data),
    .io_covSum(o_data_io_covSum)
  );
  assign io_in_a_ready = (idle | ~io_in_a_first) & i_data_ready; // @[Broadcast.scala 485:45]
  assign io_out_a_valid = o_data_io_deq_valid; // @[Broadcast.scala 496:34]
  assign io_out_a_bits_opcode = acquire ? 3'h4 : opcode; // @[Broadcast.scala 497:31]
  assign io_out_a_bits_size = size; // @[Broadcast.scala 499:25]
  assign io_out_a_bits_source = {_io_out_a_bits_source_T,source}; // @[Cat.scala 31:58]
  assign io_out_a_bits_address = address; // @[Broadcast.scala 501:25]
  assign io_out_a_bits_user_amba_prot_bufferable = user_amba_prot_bufferable; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_modifiable = user_amba_prot_modifiable; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_readalloc = user_amba_prot_readalloc; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_writealloc = user_amba_prot_writealloc; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_privileged = user_amba_prot_privileged; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_secure = user_amba_prot_secure; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_fetch = user_amba_prot_fetch; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_mask = o_data_io_deq_bits_mask; // @[Broadcast.scala 502:25]
  assign io_out_a_bits_data = o_data_io_deq_bits_data; // @[Broadcast.scala 503:25]
  assign io_source = source; // @[Broadcast.scala 478:13]
  assign io_line = address[31:6]; // @[Broadcast.scala 479:22]
  assign io_idle = got_e & sent_d; // @[Broadcast.scala 435:23]
  assign io_need_d = ~sent_d; // @[Broadcast.scala 477:16]
  assign o_data_clock = clock;
  assign o_data_reset = reset;
  assign o_data_io_enq_valid = _io_in_a_ready_T_1 & io_in_a_valid; // @[Broadcast.scala 486:44]
  assign o_data_io_enq_bits_mask = io_in_a_bits_mask; // @[Broadcast.scala 482:20 487:20]
  assign o_data_io_enq_bits_data = io_in_a_bits_data; // @[Broadcast.scala 482:20 488:20]
  assign o_data_io_deq_ready = io_out_a_ready; // @[Broadcast.scala 495:34]
  assign TLBroadcastTracker_1_covSum = 30'h0;
  assign o_data_sum = TLBroadcastTracker_1_covSum + o_data_io_covSum;
  assign io_covSum = o_data_sum;
  always @(posedge clock) begin
    got_e <= reset | _GEN_2; // @[Broadcast.scala 423:{24,24}]
    sent_d <= reset | _GEN_18; // @[Broadcast.scala 424:{24,24}]
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      opcode <= io_in_a_bits_opcode; // @[Broadcast.scala 442:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      size <= io_in_a_bits_size; // @[Broadcast.scala 444:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      source <= io_in_a_bits_source; // @[Broadcast.scala 445:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_bufferable <= io_in_a_bits_user_amba_prot_bufferable; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_modifiable <= io_in_a_bits_user_amba_prot_modifiable; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_readalloc <= io_in_a_bits_user_amba_prot_readalloc; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_writealloc <= io_in_a_bits_user_amba_prot_writealloc; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_privileged <= io_in_a_bits_user_amba_prot_privileged; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_secure <= io_in_a_bits_user_amba_prot_secure; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_fetch <= io_in_a_bits_user_amba_prot_fetch; // @[BundleMap.scala 247:19]
    end
    if (reset) begin // @[Broadcast.scala 432:24]
      address <= 32'h40; // @[Broadcast.scala 432:24]
    end else if (_T & io_in_a_first) begin
      address <= io_in_a_bits_address;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~idle & (_T_1 & ~reset)) begin
          $fatal; // @[Broadcast.scala 438:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset & ~idle) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:438 assert (idle)\n"); // @[Broadcast.scala 438:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~sent_d) & (io_d_last & _T_3)) begin
          $fatal; // @[Broadcast.scala 459:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_d_last & _T_3 & ~(~sent_d)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:459 assert (!sent_d)\n"); // @[Broadcast.scala 459:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h0 & (io_probedack & _T_3)) begin
          $fatal; // @[Broadcast.scala 468:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_probedack & _T_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:468 assert (count > 0.U)\n"); // @[Broadcast.scala 468:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  got_e = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sent_d = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  opcode = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  user_amba_prot_bufferable = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  user_amba_prot_modifiable = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  user_amba_prot_readalloc = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  user_amba_prot_writealloc = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  user_amba_prot_privileged = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  user_amba_prot_secure = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  user_amba_prot_fetch = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  address = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBroadcastTracker_2(
  input         clock,
  input         reset,
  input         io_in_a_first,
  output        io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input         io_in_a_bits_user_amba_prot_bufferable,
  input         io_in_a_bits_user_amba_prot_modifiable,
  input         io_in_a_bits_user_amba_prot_readalloc,
  input         io_in_a_bits_user_amba_prot_writealloc,
  input         io_in_a_bits_user_amba_prot_privileged,
  input         io_in_a_bits_user_amba_prot_secure,
  input         io_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  io_in_a_bits_mask,
  input  [63:0] io_in_a_bits_data,
  input         io_out_a_ready,
  output        io_out_a_valid,
  output [2:0]  io_out_a_bits_opcode,
  output [2:0]  io_out_a_bits_size,
  output [8:0]  io_out_a_bits_source,
  output [31:0] io_out_a_bits_address,
  output        io_out_a_bits_user_amba_prot_bufferable,
  output        io_out_a_bits_user_amba_prot_modifiable,
  output        io_out_a_bits_user_amba_prot_readalloc,
  output        io_out_a_bits_user_amba_prot_writealloc,
  output        io_out_a_bits_user_amba_prot_privileged,
  output        io_out_a_bits_user_amba_prot_secure,
  output        io_out_a_bits_user_amba_prot_fetch,
  output [7:0]  io_out_a_bits_mask,
  output [63:0] io_out_a_bits_data,
  input         io_probedack,
  input         io_d_last,
  output [6:0]  io_source,
  output [25:0] io_line,
  output        io_idle,
  output        io_need_d,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  o_data_clock; // @[Decoupled.scala 361:21]
  wire  o_data_reset; // @[Decoupled.scala 361:21]
  wire  o_data_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  o_data_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [7:0] o_data_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] o_data_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  o_data_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  o_data_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [7:0] o_data_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] o_data_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [29:0] o_data_io_covSum; // @[Decoupled.scala 361:21]
  reg  got_e; // @[Broadcast.scala 423:24]
  reg  sent_d; // @[Broadcast.scala 424:24]
  reg [2:0] opcode; // @[Broadcast.scala 426:20]
  reg [2:0] size; // @[Broadcast.scala 428:20]
  reg [6:0] source; // @[Broadcast.scala 429:20]
  reg  user_amba_prot_bufferable; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_modifiable; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_readalloc; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_writealloc; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_privileged; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_secure; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_fetch; // @[Broadcast.scala 430:20]
  reg [31:0] address; // @[Broadcast.scala 432:24]
  wire  idle = got_e & sent_d; // @[Broadcast.scala 435:23]
  wire  _T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = _T & io_in_a_first; // @[Broadcast.scala 437:24]
  wire  _T_3 = ~reset; // @[Broadcast.scala 438:12]
  wire  _GEN_0 = _T & io_in_a_first ? 1'h0 : sent_d; // @[Broadcast.scala 437:42 439:13 424:24]
  wire  _GEN_2 = _T & io_in_a_first ? io_in_a_bits_opcode != 3'h6 & io_in_a_bits_opcode != 3'h7 : got_e; // @[Broadcast.scala 437:42 441:13 423:24]
  wire  _GEN_18 = io_d_last | _GEN_0; // @[Broadcast.scala 458:20 460:12]
  wire  _io_in_a_ready_T_1 = idle | ~io_in_a_first; // @[Broadcast.scala 485:26]
  wire  i_data_ready = o_data_io_enq_ready; // @[Broadcast.scala 482:20 Decoupled.scala 365:17]
  wire  acquire = opcode == 3'h6 | opcode == 3'h7; // @[Broadcast.scala 491:52]
  wire [1:0] _io_out_a_bits_source_T = acquire ? 2'h3 : 2'h0; // @[Broadcast.scala 500:35]
  wire [29:0] TLBroadcastTracker_2_covSum;
  wire [29:0] o_data_sum;
  Queue_20 o_data ( // @[Decoupled.scala 361:21]
    .clock(o_data_clock),
    .reset(o_data_reset),
    .io_enq_ready(o_data_io_enq_ready),
    .io_enq_valid(o_data_io_enq_valid),
    .io_enq_bits_mask(o_data_io_enq_bits_mask),
    .io_enq_bits_data(o_data_io_enq_bits_data),
    .io_deq_ready(o_data_io_deq_ready),
    .io_deq_valid(o_data_io_deq_valid),
    .io_deq_bits_mask(o_data_io_deq_bits_mask),
    .io_deq_bits_data(o_data_io_deq_bits_data),
    .io_covSum(o_data_io_covSum)
  );
  assign io_in_a_ready = (idle | ~io_in_a_first) & i_data_ready; // @[Broadcast.scala 485:45]
  assign io_out_a_valid = o_data_io_deq_valid; // @[Broadcast.scala 496:34]
  assign io_out_a_bits_opcode = acquire ? 3'h4 : opcode; // @[Broadcast.scala 497:31]
  assign io_out_a_bits_size = size; // @[Broadcast.scala 499:25]
  assign io_out_a_bits_source = {_io_out_a_bits_source_T,source}; // @[Cat.scala 31:58]
  assign io_out_a_bits_address = address; // @[Broadcast.scala 501:25]
  assign io_out_a_bits_user_amba_prot_bufferable = user_amba_prot_bufferable; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_modifiable = user_amba_prot_modifiable; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_readalloc = user_amba_prot_readalloc; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_writealloc = user_amba_prot_writealloc; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_privileged = user_amba_prot_privileged; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_secure = user_amba_prot_secure; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_fetch = user_amba_prot_fetch; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_mask = o_data_io_deq_bits_mask; // @[Broadcast.scala 502:25]
  assign io_out_a_bits_data = o_data_io_deq_bits_data; // @[Broadcast.scala 503:25]
  assign io_source = source; // @[Broadcast.scala 478:13]
  assign io_line = address[31:6]; // @[Broadcast.scala 479:22]
  assign io_idle = got_e & sent_d; // @[Broadcast.scala 435:23]
  assign io_need_d = ~sent_d; // @[Broadcast.scala 477:16]
  assign o_data_clock = clock;
  assign o_data_reset = reset;
  assign o_data_io_enq_valid = _io_in_a_ready_T_1 & io_in_a_valid; // @[Broadcast.scala 486:44]
  assign o_data_io_enq_bits_mask = io_in_a_bits_mask; // @[Broadcast.scala 482:20 487:20]
  assign o_data_io_enq_bits_data = io_in_a_bits_data; // @[Broadcast.scala 482:20 488:20]
  assign o_data_io_deq_ready = io_out_a_ready; // @[Broadcast.scala 495:34]
  assign TLBroadcastTracker_2_covSum = 30'h0;
  assign o_data_sum = TLBroadcastTracker_2_covSum + o_data_io_covSum;
  assign io_covSum = o_data_sum;
  always @(posedge clock) begin
    got_e <= reset | _GEN_2; // @[Broadcast.scala 423:{24,24}]
    sent_d <= reset | _GEN_18; // @[Broadcast.scala 424:{24,24}]
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      opcode <= io_in_a_bits_opcode; // @[Broadcast.scala 442:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      size <= io_in_a_bits_size; // @[Broadcast.scala 444:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      source <= io_in_a_bits_source; // @[Broadcast.scala 445:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_bufferable <= io_in_a_bits_user_amba_prot_bufferable; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_modifiable <= io_in_a_bits_user_amba_prot_modifiable; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_readalloc <= io_in_a_bits_user_amba_prot_readalloc; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_writealloc <= io_in_a_bits_user_amba_prot_writealloc; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_privileged <= io_in_a_bits_user_amba_prot_privileged; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_secure <= io_in_a_bits_user_amba_prot_secure; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_fetch <= io_in_a_bits_user_amba_prot_fetch; // @[BundleMap.scala 247:19]
    end
    if (reset) begin // @[Broadcast.scala 432:24]
      address <= 32'h80; // @[Broadcast.scala 432:24]
    end else if (_T & io_in_a_first) begin
      address <= io_in_a_bits_address;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~idle & (_T_1 & ~reset)) begin
          $fatal; // @[Broadcast.scala 438:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset & ~idle) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:438 assert (idle)\n"); // @[Broadcast.scala 438:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~sent_d) & (io_d_last & _T_3)) begin
          $fatal; // @[Broadcast.scala 459:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_d_last & _T_3 & ~(~sent_d)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:459 assert (!sent_d)\n"); // @[Broadcast.scala 459:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h0 & (io_probedack & _T_3)) begin
          $fatal; // @[Broadcast.scala 468:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_probedack & _T_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:468 assert (count > 0.U)\n"); // @[Broadcast.scala 468:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  got_e = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sent_d = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  opcode = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  user_amba_prot_bufferable = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  user_amba_prot_modifiable = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  user_amba_prot_readalloc = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  user_amba_prot_writealloc = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  user_amba_prot_privileged = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  user_amba_prot_secure = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  user_amba_prot_fetch = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  address = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBroadcastTracker_3(
  input         clock,
  input         reset,
  input         io_in_a_first,
  output        io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_size,
  input  [6:0]  io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input         io_in_a_bits_user_amba_prot_bufferable,
  input         io_in_a_bits_user_amba_prot_modifiable,
  input         io_in_a_bits_user_amba_prot_readalloc,
  input         io_in_a_bits_user_amba_prot_writealloc,
  input         io_in_a_bits_user_amba_prot_privileged,
  input         io_in_a_bits_user_amba_prot_secure,
  input         io_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  io_in_a_bits_mask,
  input  [63:0] io_in_a_bits_data,
  input         io_out_a_ready,
  output        io_out_a_valid,
  output [2:0]  io_out_a_bits_opcode,
  output [2:0]  io_out_a_bits_size,
  output [8:0]  io_out_a_bits_source,
  output [31:0] io_out_a_bits_address,
  output        io_out_a_bits_user_amba_prot_bufferable,
  output        io_out_a_bits_user_amba_prot_modifiable,
  output        io_out_a_bits_user_amba_prot_readalloc,
  output        io_out_a_bits_user_amba_prot_writealloc,
  output        io_out_a_bits_user_amba_prot_privileged,
  output        io_out_a_bits_user_amba_prot_secure,
  output        io_out_a_bits_user_amba_prot_fetch,
  output [7:0]  io_out_a_bits_mask,
  output [63:0] io_out_a_bits_data,
  input         io_probedack,
  input         io_d_last,
  output [6:0]  io_source,
  output [25:0] io_line,
  output        io_idle,
  output        io_need_d,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  o_data_clock; // @[Decoupled.scala 361:21]
  wire  o_data_reset; // @[Decoupled.scala 361:21]
  wire  o_data_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  o_data_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [7:0] o_data_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] o_data_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  o_data_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  o_data_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [7:0] o_data_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] o_data_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [29:0] o_data_io_covSum; // @[Decoupled.scala 361:21]
  reg  got_e; // @[Broadcast.scala 423:24]
  reg  sent_d; // @[Broadcast.scala 424:24]
  reg [2:0] opcode; // @[Broadcast.scala 426:20]
  reg [2:0] size; // @[Broadcast.scala 428:20]
  reg [6:0] source; // @[Broadcast.scala 429:20]
  reg  user_amba_prot_bufferable; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_modifiable; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_readalloc; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_writealloc; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_privileged; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_secure; // @[Broadcast.scala 430:20]
  reg  user_amba_prot_fetch; // @[Broadcast.scala 430:20]
  reg [31:0] address; // @[Broadcast.scala 432:24]
  wire  idle = got_e & sent_d; // @[Broadcast.scala 435:23]
  wire  _T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = _T & io_in_a_first; // @[Broadcast.scala 437:24]
  wire  _T_3 = ~reset; // @[Broadcast.scala 438:12]
  wire  _GEN_0 = _T & io_in_a_first ? 1'h0 : sent_d; // @[Broadcast.scala 437:42 439:13 424:24]
  wire  _GEN_2 = _T & io_in_a_first ? io_in_a_bits_opcode != 3'h6 & io_in_a_bits_opcode != 3'h7 : got_e; // @[Broadcast.scala 437:42 441:13 423:24]
  wire  _GEN_18 = io_d_last | _GEN_0; // @[Broadcast.scala 458:20 460:12]
  wire  _io_in_a_ready_T_1 = idle | ~io_in_a_first; // @[Broadcast.scala 485:26]
  wire  i_data_ready = o_data_io_enq_ready; // @[Broadcast.scala 482:20 Decoupled.scala 365:17]
  wire  acquire = opcode == 3'h6 | opcode == 3'h7; // @[Broadcast.scala 491:52]
  wire [1:0] _io_out_a_bits_source_T = acquire ? 2'h3 : 2'h0; // @[Broadcast.scala 500:35]
  wire [29:0] TLBroadcastTracker_3_covSum;
  wire [29:0] o_data_sum;
  Queue_20 o_data ( // @[Decoupled.scala 361:21]
    .clock(o_data_clock),
    .reset(o_data_reset),
    .io_enq_ready(o_data_io_enq_ready),
    .io_enq_valid(o_data_io_enq_valid),
    .io_enq_bits_mask(o_data_io_enq_bits_mask),
    .io_enq_bits_data(o_data_io_enq_bits_data),
    .io_deq_ready(o_data_io_deq_ready),
    .io_deq_valid(o_data_io_deq_valid),
    .io_deq_bits_mask(o_data_io_deq_bits_mask),
    .io_deq_bits_data(o_data_io_deq_bits_data),
    .io_covSum(o_data_io_covSum)
  );
  assign io_in_a_ready = (idle | ~io_in_a_first) & i_data_ready; // @[Broadcast.scala 485:45]
  assign io_out_a_valid = o_data_io_deq_valid; // @[Broadcast.scala 496:34]
  assign io_out_a_bits_opcode = acquire ? 3'h4 : opcode; // @[Broadcast.scala 497:31]
  assign io_out_a_bits_size = size; // @[Broadcast.scala 499:25]
  assign io_out_a_bits_source = {_io_out_a_bits_source_T,source}; // @[Cat.scala 31:58]
  assign io_out_a_bits_address = address; // @[Broadcast.scala 501:25]
  assign io_out_a_bits_user_amba_prot_bufferable = user_amba_prot_bufferable; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_modifiable = user_amba_prot_modifiable; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_readalloc = user_amba_prot_readalloc; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_writealloc = user_amba_prot_writealloc; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_privileged = user_amba_prot_privileged; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_secure = user_amba_prot_secure; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_user_amba_prot_fetch = user_amba_prot_fetch; // @[BundleMap.scala 247:19]
  assign io_out_a_bits_mask = o_data_io_deq_bits_mask; // @[Broadcast.scala 502:25]
  assign io_out_a_bits_data = o_data_io_deq_bits_data; // @[Broadcast.scala 503:25]
  assign io_source = source; // @[Broadcast.scala 478:13]
  assign io_line = address[31:6]; // @[Broadcast.scala 479:22]
  assign io_idle = got_e & sent_d; // @[Broadcast.scala 435:23]
  assign io_need_d = ~sent_d; // @[Broadcast.scala 477:16]
  assign o_data_clock = clock;
  assign o_data_reset = reset;
  assign o_data_io_enq_valid = _io_in_a_ready_T_1 & io_in_a_valid; // @[Broadcast.scala 486:44]
  assign o_data_io_enq_bits_mask = io_in_a_bits_mask; // @[Broadcast.scala 482:20 487:20]
  assign o_data_io_enq_bits_data = io_in_a_bits_data; // @[Broadcast.scala 482:20 488:20]
  assign o_data_io_deq_ready = io_out_a_ready; // @[Broadcast.scala 495:34]
  assign TLBroadcastTracker_3_covSum = 30'h0;
  assign o_data_sum = TLBroadcastTracker_3_covSum + o_data_io_covSum;
  assign io_covSum = o_data_sum;
  always @(posedge clock) begin
    got_e <= reset | _GEN_2; // @[Broadcast.scala 423:{24,24}]
    sent_d <= reset | _GEN_18; // @[Broadcast.scala 424:{24,24}]
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      opcode <= io_in_a_bits_opcode; // @[Broadcast.scala 442:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      size <= io_in_a_bits_size; // @[Broadcast.scala 444:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      source <= io_in_a_bits_source; // @[Broadcast.scala 445:13]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_bufferable <= io_in_a_bits_user_amba_prot_bufferable; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_modifiable <= io_in_a_bits_user_amba_prot_modifiable; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_readalloc <= io_in_a_bits_user_amba_prot_readalloc; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_writealloc <= io_in_a_bits_user_amba_prot_writealloc; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_privileged <= io_in_a_bits_user_amba_prot_privileged; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_secure <= io_in_a_bits_user_amba_prot_secure; // @[BundleMap.scala 247:19]
    end
    if (_T & io_in_a_first) begin // @[Broadcast.scala 437:42]
      user_amba_prot_fetch <= io_in_a_bits_user_amba_prot_fetch; // @[BundleMap.scala 247:19]
    end
    if (reset) begin // @[Broadcast.scala 432:24]
      address <= 32'hc0; // @[Broadcast.scala 432:24]
    end else if (_T & io_in_a_first) begin
      address <= io_in_a_bits_address;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~idle & (_T_1 & ~reset)) begin
          $fatal; // @[Broadcast.scala 438:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset & ~idle) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:438 assert (idle)\n"); // @[Broadcast.scala 438:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~sent_d) & (io_d_last & _T_3)) begin
          $fatal; // @[Broadcast.scala 459:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_d_last & _T_3 & ~(~sent_d)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:459 assert (!sent_d)\n"); // @[Broadcast.scala 459:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h0 & (io_probedack & _T_3)) begin
          $fatal; // @[Broadcast.scala 468:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_probedack & _T_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:468 assert (count > 0.U)\n"); // @[Broadcast.scala 468:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  got_e = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sent_d = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  opcode = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  user_amba_prot_bufferable = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  user_amba_prot_modifiable = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  user_amba_prot_readalloc = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  user_amba_prot_writealloc = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  user_amba_prot_privileged = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  user_amba_prot_secure = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  user_amba_prot_fetch = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  address = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBroadcast(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_size,
  input  [6:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input         auto_in_a_bits_user_amba_prot_bufferable,
  input         auto_in_a_bits_user_amba_prot_modifiable,
  input         auto_in_a_bits_user_amba_prot_readalloc,
  input         auto_in_a_bits_user_amba_prot_writealloc,
  input         auto_in_a_bits_user_amba_prot_privileged,
  input         auto_in_a_bits_user_amba_prot_secure,
  input         auto_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [2:0]  auto_in_d_bits_size,
  output [6:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_size,
  output [8:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output        auto_out_a_bits_user_amba_prot_bufferable,
  output        auto_out_a_bits_user_amba_prot_modifiable,
  output        auto_out_a_bits_user_amba_prot_readalloc,
  output        auto_out_a_bits_user_amba_prot_writealloc,
  output        auto_out_a_bits_user_amba_prot_privileged,
  output        auto_out_a_bits_user_amba_prot_secure,
  output        auto_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [2:0]  auto_out_d_bits_size,
  input  [8:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  BroadcastFilter_io_request_ready; // @[Broadcast.scala 99:26]
  wire  BroadcastFilter_io_request_valid; // @[Broadcast.scala 99:26]
  wire  BroadcastFilter_io_response_ready; // @[Broadcast.scala 99:26]
  wire  BroadcastFilter_io_response_valid; // @[Broadcast.scala 99:26]
  wire [29:0] BroadcastFilter_io_covSum; // @[Broadcast.scala 99:26]
  wire  TLBroadcastTracker_clock; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_reset; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_first; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_ready; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_valid; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_io_in_a_bits_opcode; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_io_in_a_bits_size; // @[Broadcast.scala 107:15]
  wire [6:0] TLBroadcastTracker_io_in_a_bits_source; // @[Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_io_in_a_bits_address; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_bits_user_amba_prot_bufferable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_bits_user_amba_prot_modifiable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_bits_user_amba_prot_readalloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_bits_user_amba_prot_writealloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_bits_user_amba_prot_privileged; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_bits_user_amba_prot_secure; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_bits_user_amba_prot_fetch; // @[Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_io_in_a_bits_mask; // @[Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_io_in_a_bits_data; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_ready; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_valid; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_io_out_a_bits_opcode; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_io_out_a_bits_size; // @[Broadcast.scala 107:15]
  wire [8:0] TLBroadcastTracker_io_out_a_bits_source; // @[Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_io_out_a_bits_address; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_bits_user_amba_prot_bufferable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_bits_user_amba_prot_modifiable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_bits_user_amba_prot_readalloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_bits_user_amba_prot_writealloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_bits_user_amba_prot_privileged; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_bits_user_amba_prot_secure; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_bits_user_amba_prot_fetch; // @[Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_io_out_a_bits_mask; // @[Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_io_out_a_bits_data; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_probedack; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_d_last; // @[Broadcast.scala 107:15]
  wire [6:0] TLBroadcastTracker_io_source; // @[Broadcast.scala 107:15]
  wire [25:0] TLBroadcastTracker_io_line; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_idle; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_need_d; // @[Broadcast.scala 107:15]
  wire [29:0] TLBroadcastTracker_io_covSum; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_clock; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_reset; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_first; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_ready; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_valid; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_1_io_in_a_bits_opcode; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_1_io_in_a_bits_size; // @[Broadcast.scala 107:15]
  wire [6:0] TLBroadcastTracker_1_io_in_a_bits_source; // @[Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_1_io_in_a_bits_address; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_bufferable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_modifiable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_readalloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_writealloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_privileged; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_secure; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_fetch; // @[Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_1_io_in_a_bits_mask; // @[Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_1_io_in_a_bits_data; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_ready; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_valid; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_1_io_out_a_bits_opcode; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_1_io_out_a_bits_size; // @[Broadcast.scala 107:15]
  wire [8:0] TLBroadcastTracker_1_io_out_a_bits_source; // @[Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_1_io_out_a_bits_address; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_bufferable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_modifiable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_readalloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_writealloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_privileged; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_secure; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_fetch; // @[Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_1_io_out_a_bits_mask; // @[Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_1_io_out_a_bits_data; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_probedack; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_d_last; // @[Broadcast.scala 107:15]
  wire [6:0] TLBroadcastTracker_1_io_source; // @[Broadcast.scala 107:15]
  wire [25:0] TLBroadcastTracker_1_io_line; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_idle; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_need_d; // @[Broadcast.scala 107:15]
  wire [29:0] TLBroadcastTracker_1_io_covSum; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_clock; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_reset; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_first; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_ready; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_valid; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_2_io_in_a_bits_opcode; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_2_io_in_a_bits_size; // @[Broadcast.scala 107:15]
  wire [6:0] TLBroadcastTracker_2_io_in_a_bits_source; // @[Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_2_io_in_a_bits_address; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_bufferable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_modifiable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_readalloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_writealloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_privileged; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_secure; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_fetch; // @[Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_2_io_in_a_bits_mask; // @[Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_2_io_in_a_bits_data; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_ready; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_valid; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_2_io_out_a_bits_opcode; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_2_io_out_a_bits_size; // @[Broadcast.scala 107:15]
  wire [8:0] TLBroadcastTracker_2_io_out_a_bits_source; // @[Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_2_io_out_a_bits_address; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_bufferable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_modifiable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_readalloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_writealloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_privileged; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_secure; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_fetch; // @[Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_2_io_out_a_bits_mask; // @[Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_2_io_out_a_bits_data; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_probedack; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_d_last; // @[Broadcast.scala 107:15]
  wire [6:0] TLBroadcastTracker_2_io_source; // @[Broadcast.scala 107:15]
  wire [25:0] TLBroadcastTracker_2_io_line; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_idle; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_need_d; // @[Broadcast.scala 107:15]
  wire [29:0] TLBroadcastTracker_2_io_covSum; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_clock; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_reset; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_first; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_ready; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_valid; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_3_io_in_a_bits_opcode; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_3_io_in_a_bits_size; // @[Broadcast.scala 107:15]
  wire [6:0] TLBroadcastTracker_3_io_in_a_bits_source; // @[Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_3_io_in_a_bits_address; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_bufferable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_modifiable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_readalloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_writealloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_privileged; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_secure; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_fetch; // @[Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_3_io_in_a_bits_mask; // @[Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_3_io_in_a_bits_data; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_ready; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_valid; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_3_io_out_a_bits_opcode; // @[Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_3_io_out_a_bits_size; // @[Broadcast.scala 107:15]
  wire [8:0] TLBroadcastTracker_3_io_out_a_bits_source; // @[Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_3_io_out_a_bits_address; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_bufferable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_modifiable; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_readalloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_writealloc; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_privileged; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_secure; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_fetch; // @[Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_3_io_out_a_bits_mask; // @[Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_3_io_out_a_bits_data; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_probedack; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_d_last; // @[Broadcast.scala 107:15]
  wire [6:0] TLBroadcastTracker_3_io_source; // @[Broadcast.scala 107:15]
  wire [25:0] TLBroadcastTracker_3_io_line; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_idle; // @[Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_need_d; // @[Broadcast.scala 107:15]
  wire [29:0] TLBroadcastTracker_3_io_covSum; // @[Broadcast.scala 107:15]
  wire  _T_14 = auto_out_d_bits_source[8:7] == 2'h1; // @[Broadcast.scala 119:27]
  wire  opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [2:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 3'h0; // @[Arbiter.scala 88:28]
  wire  _T_56 = opdata | ~auto_out_d_bits_source[8]; // @[Broadcast.scala 140:34]
  reg [2:0] counter; // @[Edges.scala 228:27]
  wire [2:0] _T_38 = opdata ? 3'h5 : 3'h6; // @[Broadcast.scala 132:36]
  wire [2:0] out_1_bits_opcode = auto_out_d_bits_source[8] ? _T_38 : auto_out_d_bits_opcode; // @[Broadcast.scala 130:21 131:24 132:30]
  wire  beats1_opdata = out_1_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [12:0] _beats1_decode_T_1 = 13'h3f << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire [2:0] beats1_decode = _beats1_decode_T_3[5:3]; // @[Edges.scala 219:59]
  wire [2:0] beats1 = beats1_opdata ? beats1_decode : 3'h0; // @[Edges.scala 220:14]
  wire  last = counter == 3'h1 | beats1 == 3'h0; // @[Edges.scala 231:37]
  wire  _T_35 = ~_T_14; // @[Broadcast.scala 129:51]
  wire  out_1_earlyValid = auto_out_d_valid & ~_T_14; // @[Broadcast.scala 129:48]
  wire [1:0] _readys_T = {out_1_earlyValid,1'h0}; // @[Cat.scala 31:58]
  wire [2:0] _readys_T_1 = {_readys_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0]; // @[package.scala 244:43]
  wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0}; // @[Arbiter.scala 16:78]
  wire [1:0] _readys_T_7 = ~_readys_T_5[1:0]; // @[Arbiter.scala 16:61]
  wire  readys__1 = _readys_T_7[1]; // @[Arbiter.scala 95:86]
  reg  state__1; // @[Arbiter.scala 116:26]
  wire  allowed__1 = idle ? readys__1 : state__1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_in_d_ready & allowed__1; // @[Arbiter.scala 123:31]
  wire  _T_15 = out_1_ready & out_1_earlyValid; // @[Decoupled.scala 50:35]
  wire [2:0] counter1 = counter - 3'h1; // @[Edges.scala 229:28]
  wire  first = counter == 3'h0; // @[Edges.scala 230:25]
  wire [6:0] out_1_bits_source = auto_out_d_bits_source[6:0]; // @[Broadcast.scala 121:26 130:21]
  wire  _T_17 = TLBroadcastTracker_io_need_d & TLBroadcastTracker_io_source == out_1_bits_source; // @[Broadcast.scala 123:62]
  wire  _T_19 = TLBroadcastTracker_1_io_need_d & TLBroadcastTracker_1_io_source == out_1_bits_source; // @[Broadcast.scala 123:62]
  wire  _T_21 = TLBroadcastTracker_2_io_need_d & TLBroadcastTracker_2_io_source == out_1_bits_source; // @[Broadcast.scala 123:62]
  wire  _T_23 = TLBroadcastTracker_3_io_need_d & TLBroadcastTracker_3_io_source == out_1_bits_source; // @[Broadcast.scala 123:62]
  wire [3:0] _T_24 = {_T_23,_T_21,_T_19,_T_17}; // @[Broadcast.scala 123:102]
  reg [3:0] r; // @[Reg.scala 16:16]
  wire [3:0] _GEN_1 = first ? _T_24 : r; // @[Reg.scala 16:16 17:{18,22}]
  wire  _T_32 = ~reset; // @[Broadcast.scala 125:14]
  wire  bundleOut_0_d_ready = out_1_ready | _T_14; // @[Broadcast.scala 128:50]
  wire  _T_46 = ~out_1_earlyValid; // @[Broadcast.scala 137:15]
  wire  _T_65 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  reg [2:0] beatsLeft_1; // @[Arbiter.scala 87:30]
  wire  idle_1 = beatsLeft_1 == 3'h0; // @[Arbiter.scala 88:28]
  wire  out_7_earlyValid = TLBroadcastTracker_3_io_out_a_valid; // @[ReadyValidCancel.scala 68:19 69:20]
  wire  out_6_earlyValid = TLBroadcastTracker_2_io_out_a_valid; // @[ReadyValidCancel.scala 68:19 69:20]
  wire  out_5_earlyValid = TLBroadcastTracker_1_io_out_a_valid; // @[ReadyValidCancel.scala 68:19 69:20]
  wire  out_4_earlyValid = TLBroadcastTracker_io_out_a_valid; // @[ReadyValidCancel.scala 68:19 69:20]
  wire [4:0] _readys_T_10 = {out_7_earlyValid,out_6_earlyValid,out_5_earlyValid,out_4_earlyValid,1'h0}; // @[Cat.scala 31:58]
  wire [5:0] _readys_T_11 = {_readys_T_10, 1'h0}; // @[package.scala 244:48]
  wire [4:0] _readys_T_13 = _readys_T_10 | _readys_T_11[4:0]; // @[package.scala 244:43]
  wire [6:0] _readys_T_14 = {_readys_T_13, 2'h0}; // @[package.scala 244:48]
  wire [4:0] _readys_T_16 = _readys_T_13 | _readys_T_14[4:0]; // @[package.scala 244:43]
  wire [8:0] _readys_T_17 = {_readys_T_16, 4'h0}; // @[package.scala 244:48]
  wire [4:0] _readys_T_19 = _readys_T_16 | _readys_T_17[4:0]; // @[package.scala 244:43]
  wire [5:0] _readys_T_21 = {_readys_T_19, 1'h0}; // @[Arbiter.scala 16:78]
  wire [4:0] _readys_T_23 = ~_readys_T_21[4:0]; // @[Arbiter.scala 16:61]
  wire  latch = idle & auto_in_d_ready; // @[Arbiter.scala 89:24]
  wire  earlyWinner__1 = readys__1 & out_1_earlyValid; // @[Arbiter.scala 97:79]
  wire  muxStateEarly__1 = idle ? earlyWinner__1 : state__1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_2 = state__1 & out_1_earlyValid; // @[Mux.scala 27:73]
  wire  sink_ACancel_earlyValid = idle ? out_1_earlyValid : _sink_ACancel_earlyValid_T_2; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_in_d_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [2:0] _GEN_3 = {{2'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [2:0] _beatsLeft_T_4 = beatsLeft - _GEN_3; // @[Arbiter.scala 113:52]
  wire [12:0] _decode_T_13 = 13'h3f << TLBroadcastTracker_io_out_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _decode_T_15 = ~_decode_T_13[5:0]; // @[package.scala 234:46]
  wire [2:0] decode_3 = _decode_T_15[5:3]; // @[Edges.scala 219:59]
  wire  opdata_4 = ~TLBroadcastTracker_io_out_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [2:0] _T_257 = opdata_4 ? decode_3 : 3'h0; // @[Edges.scala 220:14]
  wire [12:0] _decode_T_17 = 13'h3f << TLBroadcastTracker_1_io_out_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _decode_T_19 = ~_decode_T_17[5:0]; // @[package.scala 234:46]
  wire [2:0] decode_4 = _decode_T_19[5:3]; // @[Edges.scala 219:59]
  wire  opdata_5 = ~TLBroadcastTracker_1_io_out_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [2:0] _T_258 = opdata_5 ? decode_4 : 3'h0; // @[Edges.scala 220:14]
  wire [12:0] _decode_T_21 = 13'h3f << TLBroadcastTracker_2_io_out_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _decode_T_23 = ~_decode_T_21[5:0]; // @[package.scala 234:46]
  wire [2:0] decode_5 = _decode_T_23[5:3]; // @[Edges.scala 219:59]
  wire  opdata_6 = ~TLBroadcastTracker_2_io_out_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [2:0] _T_259 = opdata_6 ? decode_5 : 3'h0; // @[Edges.scala 220:14]
  wire [12:0] _decode_T_25 = 13'h3f << TLBroadcastTracker_3_io_out_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _decode_T_27 = ~_decode_T_25[5:0]; // @[package.scala 234:46]
  wire [2:0] decode_6 = _decode_T_27[5:3]; // @[Edges.scala 219:59]
  wire  opdata_7 = ~TLBroadcastTracker_3_io_out_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [2:0] _T_260 = opdata_7 ? decode_6 : 3'h0; // @[Edges.scala 220:14]
  wire  latch_1 = idle_1 & auto_out_a_ready; // @[Arbiter.scala 89:24]
  wire  readys_1_1 = _readys_T_23[1]; // @[Arbiter.scala 95:86]
  wire  readys_1_2 = _readys_T_23[2]; // @[Arbiter.scala 95:86]
  wire  readys_1_3 = _readys_T_23[3]; // @[Arbiter.scala 95:86]
  wire  readys_1_4 = _readys_T_23[4]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_1_1 = readys_1_1 & out_4_earlyValid; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1_2 = readys_1_2 & out_5_earlyValid; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1_3 = readys_1_3 & out_6_earlyValid; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1_4 = readys_1_4 & out_7_earlyValid; // @[Arbiter.scala 97:79]
  wire  prefixOR_3 = earlyWinner_1_1 | earlyWinner_1_2; // @[Arbiter.scala 104:53]
  wire  prefixOR_4 = prefixOR_3 | earlyWinner_1_3; // @[Arbiter.scala 104:53]
  wire  _T_286 = out_4_earlyValid | out_5_earlyValid | out_6_earlyValid | out_7_earlyValid; // @[Arbiter.scala 107:36]
  wire  _T_287 = ~(out_4_earlyValid | out_5_earlyValid | out_6_earlyValid | out_7_earlyValid); // @[Arbiter.scala 107:15]
  wire [2:0] maskedBeats_1_1 = earlyWinner_1_1 ? _T_257 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_2 = earlyWinner_1_2 ? _T_258 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_3 = earlyWinner_1_3 ? _T_259 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] maskedBeats_4 = earlyWinner_1_4 ? _T_260 : 3'h0; // @[Arbiter.scala 111:73]
  wire [2:0] _initBeats_T_1 = maskedBeats_1_1 | maskedBeats_2; // @[Arbiter.scala 112:44]
  wire [2:0] _initBeats_T_2 = _initBeats_T_1 | maskedBeats_3; // @[Arbiter.scala 112:44]
  wire [2:0] initBeats_1 = _initBeats_T_2 | maskedBeats_4; // @[Arbiter.scala 112:44]
  reg  state_1_1; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_1_1 = idle_1 ? earlyWinner_1_1 : state_1_1; // @[Arbiter.scala 117:30]
  reg  state_1_2; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_1_2 = idle_1 ? earlyWinner_1_2 : state_1_2; // @[Arbiter.scala 117:30]
  reg  state_1_3; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_1_3 = idle_1 ? earlyWinner_1_3 : state_1_3; // @[Arbiter.scala 117:30]
  reg  state_1_4; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_1_4 = idle_1 ? earlyWinner_1_4 : state_1_4; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_17 = state_1_1 & out_4_earlyValid | state_1_2 & out_5_earlyValid | state_1_3 &
    out_6_earlyValid | state_1_4 & out_7_earlyValid; // @[Mux.scala 27:73]
  wire  sink_ACancel_1_earlyValid = idle_1 ? _T_286 : _sink_ACancel_earlyValid_T_17; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_8 = auto_out_a_ready & sink_ACancel_1_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [2:0] _GEN_8 = {{2'd0}, _beatsLeft_T_8}; // @[Arbiter.scala 113:52]
  wire [2:0] _beatsLeft_T_10 = beatsLeft_1 - _GEN_8; // @[Arbiter.scala 113:52]
  wire  allowed_1_1 = idle_1 ? readys_1_1 : state_1_1; // @[Arbiter.scala 121:24]
  wire  allowed_1_2 = idle_1 ? readys_1_2 : state_1_2; // @[Arbiter.scala 121:24]
  wire  allowed_1_3 = idle_1 ? readys_1_3 : state_1_3; // @[Arbiter.scala 121:24]
  wire  allowed_1_4 = idle_1 ? readys_1_4 : state_1_4; // @[Arbiter.scala 121:24]
  wire [63:0] out_4_bits_data = TLBroadcastTracker_io_out_a_bits_data; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [63:0] _T_319 = muxStateEarly_1_1 ? out_4_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] out_5_bits_data = TLBroadcastTracker_1_io_out_a_bits_data; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [63:0] _T_320 = muxStateEarly_1_2 ? out_5_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] out_6_bits_data = TLBroadcastTracker_2_io_out_a_bits_data; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [63:0] _T_321 = muxStateEarly_1_3 ? out_6_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] out_7_bits_data = TLBroadcastTracker_3_io_out_a_bits_data; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [63:0] _T_322 = muxStateEarly_1_4 ? out_7_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_324 = _T_319 | _T_320; // @[Mux.scala 27:73]
  wire [63:0] _T_325 = _T_324 | _T_321; // @[Mux.scala 27:73]
  wire [7:0] out_4_bits_mask = TLBroadcastTracker_io_out_a_bits_mask; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [7:0] _T_328 = muxStateEarly_1_1 ? out_4_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] out_5_bits_mask = TLBroadcastTracker_1_io_out_a_bits_mask; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [7:0] _T_329 = muxStateEarly_1_2 ? out_5_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] out_6_bits_mask = TLBroadcastTracker_2_io_out_a_bits_mask; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [7:0] _T_330 = muxStateEarly_1_3 ? out_6_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] out_7_bits_mask = TLBroadcastTracker_3_io_out_a_bits_mask; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [7:0] _T_331 = muxStateEarly_1_4 ? out_7_bits_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_333 = _T_328 | _T_329; // @[Mux.scala 27:73]
  wire [7:0] _T_334 = _T_333 | _T_330; // @[Mux.scala 27:73]
  wire  out_4_bits_user_amba_prot_fetch = TLBroadcastTracker_io_out_a_bits_user_amba_prot_fetch; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_5_bits_user_amba_prot_fetch = TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_fetch; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_6_bits_user_amba_prot_fetch = TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_fetch; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_7_bits_user_amba_prot_fetch = TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_fetch; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_4_bits_user_amba_prot_secure = TLBroadcastTracker_io_out_a_bits_user_amba_prot_secure; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_5_bits_user_amba_prot_secure = TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_secure; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_6_bits_user_amba_prot_secure = TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_secure; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_7_bits_user_amba_prot_secure = TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_secure; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_4_bits_user_amba_prot_privileged = TLBroadcastTracker_io_out_a_bits_user_amba_prot_privileged; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_5_bits_user_amba_prot_privileged = TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_privileged; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_6_bits_user_amba_prot_privileged = TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_privileged; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_7_bits_user_amba_prot_privileged = TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_privileged; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_4_bits_user_amba_prot_writealloc = TLBroadcastTracker_io_out_a_bits_user_amba_prot_writealloc; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_5_bits_user_amba_prot_writealloc = TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_writealloc; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_6_bits_user_amba_prot_writealloc = TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_writealloc; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_7_bits_user_amba_prot_writealloc = TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_writealloc; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_4_bits_user_amba_prot_readalloc = TLBroadcastTracker_io_out_a_bits_user_amba_prot_readalloc; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_5_bits_user_amba_prot_readalloc = TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_readalloc; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_6_bits_user_amba_prot_readalloc = TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_readalloc; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_7_bits_user_amba_prot_readalloc = TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_readalloc; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_4_bits_user_amba_prot_modifiable = TLBroadcastTracker_io_out_a_bits_user_amba_prot_modifiable; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_5_bits_user_amba_prot_modifiable = TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_modifiable; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_6_bits_user_amba_prot_modifiable = TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_modifiable; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_7_bits_user_amba_prot_modifiable = TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_modifiable; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_4_bits_user_amba_prot_bufferable = TLBroadcastTracker_io_out_a_bits_user_amba_prot_bufferable; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_5_bits_user_amba_prot_bufferable = TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_bufferable; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_6_bits_user_amba_prot_bufferable = TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_bufferable; // @[ReadyValidCancel.scala 68:19 71:14]
  wire  out_7_bits_user_amba_prot_bufferable = TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_bufferable; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [31:0] out_4_bits_address = TLBroadcastTracker_io_out_a_bits_address; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [31:0] _T_400 = muxStateEarly_1_1 ? out_4_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] out_5_bits_address = TLBroadcastTracker_1_io_out_a_bits_address; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [31:0] _T_401 = muxStateEarly_1_2 ? out_5_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] out_6_bits_address = TLBroadcastTracker_2_io_out_a_bits_address; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [31:0] _T_402 = muxStateEarly_1_3 ? out_6_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] out_7_bits_address = TLBroadcastTracker_3_io_out_a_bits_address; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [31:0] _T_403 = muxStateEarly_1_4 ? out_7_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_405 = _T_400 | _T_401; // @[Mux.scala 27:73]
  wire [31:0] _T_406 = _T_405 | _T_402; // @[Mux.scala 27:73]
  wire [8:0] out_4_bits_source = TLBroadcastTracker_io_out_a_bits_source; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [8:0] _T_409 = muxStateEarly_1_1 ? out_4_bits_source : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] out_5_bits_source = TLBroadcastTracker_1_io_out_a_bits_source; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [8:0] _T_410 = muxStateEarly_1_2 ? out_5_bits_source : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] out_6_bits_source = TLBroadcastTracker_2_io_out_a_bits_source; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [8:0] _T_411 = muxStateEarly_1_3 ? out_6_bits_source : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] out_7_bits_source = TLBroadcastTracker_3_io_out_a_bits_source; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [8:0] _T_412 = muxStateEarly_1_4 ? out_7_bits_source : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _T_414 = _T_409 | _T_410; // @[Mux.scala 27:73]
  wire [8:0] _T_415 = _T_414 | _T_411; // @[Mux.scala 27:73]
  wire [2:0] out_4_bits_size = TLBroadcastTracker_io_out_a_bits_size; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_418 = muxStateEarly_1_1 ? out_4_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] out_5_bits_size = TLBroadcastTracker_1_io_out_a_bits_size; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_419 = muxStateEarly_1_2 ? out_5_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] out_6_bits_size = TLBroadcastTracker_2_io_out_a_bits_size; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_420 = muxStateEarly_1_3 ? out_6_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] out_7_bits_size = TLBroadcastTracker_3_io_out_a_bits_size; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_421 = muxStateEarly_1_4 ? out_7_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_423 = _T_418 | _T_419; // @[Mux.scala 27:73]
  wire [2:0] _T_424 = _T_423 | _T_420; // @[Mux.scala 27:73]
  wire [2:0] out_4_bits_opcode = TLBroadcastTracker_io_out_a_bits_opcode; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_436 = muxStateEarly_1_1 ? out_4_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] out_5_bits_opcode = TLBroadcastTracker_1_io_out_a_bits_opcode; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_437 = muxStateEarly_1_2 ? out_5_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] out_6_bits_opcode = TLBroadcastTracker_2_io_out_a_bits_opcode; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_438 = muxStateEarly_1_3 ? out_6_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] out_7_bits_opcode = TLBroadcastTracker_3_io_out_a_bits_opcode; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_439 = muxStateEarly_1_4 ? out_7_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_441 = _T_436 | _T_437; // @[Mux.scala 27:73]
  wire [2:0] _T_442 = _T_441 | _T_438; // @[Mux.scala 27:73]
  reg  REG; // @[Broadcast.scala 215:31]
  wire [1:0] _GEN_9 = {{1'd0}, REG}; // @[Broadcast.scala 218:35]
  wire  _T_448 = |REG; // @[Broadcast.scala 219:38]
  reg [2:0] counter_2; // @[Edges.scala 228:27]
  wire  first_2 = counter_2 == 3'h0; // @[Edges.scala 230:25]
  wire  _bundleIn_0_a_ready_T_1 = ~first_2 | BroadcastFilter_io_request_ready; // @[Broadcast.scala 243:31]
  wire [3:0] _T_463 = {TLBroadcastTracker_3_io_line == auto_in_a_bits_address[31:6],TLBroadcastTracker_2_io_line ==
    auto_in_a_bits_address[31:6],TLBroadcastTracker_1_io_line == auto_in_a_bits_address[31:6],TLBroadcastTracker_io_line
     == auto_in_a_bits_address[31:6]}; // @[Broadcast.scala 236:100]
  wire  _T_464 = |_T_463; // @[Broadcast.scala 237:43]
  wire  _WIRE_85_3 = TLBroadcastTracker_3_io_idle; // @[Broadcast.scala 234:{33,33}]
  wire  _WIRE_85_2 = TLBroadcastTracker_2_io_idle; // @[Broadcast.scala 234:{33,33}]
  wire  _WIRE_85_1 = TLBroadcastTracker_1_io_idle; // @[Broadcast.scala 234:{33,33}]
  wire  _WIRE_85_0 = TLBroadcastTracker_io_idle; // @[Broadcast.scala 234:{33,33}]
  wire [3:0] _T_453 = {_WIRE_85_3,_WIRE_85_2,_WIRE_85_1,_WIRE_85_0}; // @[Broadcast.scala 234:64]
  wire [4:0] _T_465 = {_T_453, 1'h0}; // @[package.scala 244:48]
  wire [3:0] _T_467 = _T_453 | _T_465[3:0]; // @[package.scala 244:43]
  wire [5:0] _T_468 = {_T_467, 2'h0}; // @[package.scala 244:48]
  wire [3:0] _T_470 = _T_467 | _T_468[3:0]; // @[package.scala 244:43]
  wire [4:0] _T_472 = {_T_470, 1'h0}; // @[Broadcast.scala 238:64]
  wire [4:0] _T_473 = ~_T_472; // @[Broadcast.scala 238:41]
  wire [4:0] _GEN_15 = {{1'd0}, _T_453}; // @[Broadcast.scala 238:39]
  wire [4:0] _T_474 = _GEN_15 & _T_473; // @[Broadcast.scala 238:39]
  wire [4:0] _T_475 = _T_464 ? {{1'd0}, _T_463} : _T_474; // @[Broadcast.scala 239:30]
  wire  _WIRE_87_3 = TLBroadcastTracker_3_io_in_a_ready; // @[Broadcast.scala 240:{34,34}]
  wire  _WIRE_87_2 = TLBroadcastTracker_2_io_in_a_ready; // @[Broadcast.scala 240:{34,34}]
  wire  _WIRE_87_1 = TLBroadcastTracker_1_io_in_a_ready; // @[Broadcast.scala 240:{34,34}]
  wire  _WIRE_87_0 = TLBroadcastTracker_io_in_a_ready; // @[Broadcast.scala 240:{34,34}]
  wire [3:0] _T_476 = {_WIRE_87_3,_WIRE_87_2,_WIRE_87_1,_WIRE_87_0}; // @[Broadcast.scala 240:63]
  wire [4:0] _GEN_16 = {{1'd0}, _T_476}; // @[Broadcast.scala 241:41]
  wire [4:0] _T_477 = _T_475 & _GEN_16; // @[Broadcast.scala 241:41]
  wire  _T_478 = |_T_477; // @[Broadcast.scala 241:61]
  wire  bundleIn_0_a_ready = (~first_2 | BroadcastFilter_io_request_ready) & _T_478; // @[Broadcast.scala 243:59]
  wire  _T_452 = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 50:35]
  wire [12:0] _beats1_decode_T_9 = 13'h3f << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_11 = ~_beats1_decode_T_9[5:0]; // @[package.scala 234:46]
  wire [2:0] beats1_decode_2 = _beats1_decode_T_11[5:3]; // @[Edges.scala 219:59]
  wire  beats1_opdata_2 = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [2:0] counter1_2 = counter_2 - 3'h1; // @[Edges.scala 229:28]
  wire  _T_534 = BroadcastFilter_io_response_ready & BroadcastFilter_io_response_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_7 = _T_534 ? 2'h0 : _GEN_9; // @[Broadcast.scala 260:40 261:21]
  reg [4:0] TLBroadcast_covState; // @[Register tracking TLBroadcast state]
  reg  TLBroadcast_covMap [0:31]; // @[Coverage map for TLBroadcast]
  wire  TLBroadcast_covMap_read_en; // @[Coverage map for TLBroadcast]
  wire [4:0] TLBroadcast_covMap_read_addr; // @[Coverage map for TLBroadcast]
  wire  TLBroadcast_covMap_read_data; // @[Coverage map for TLBroadcast]
  wire  TLBroadcast_covMap_write_data; // @[Coverage map for TLBroadcast]
  wire [4:0] TLBroadcast_covMap_write_addr; // @[Coverage map for TLBroadcast]
  wire  TLBroadcast_covMap_write_mask; // @[Coverage map for TLBroadcast]
  wire  TLBroadcast_covMap_write_en; // @[Coverage map for TLBroadcast]
  reg [29:0] TLBroadcast_covSum; // @[Sum of coverage map]
  wire  state_1_3_shl;
  wire [4:0] state_1_3_pad;
  wire [1:0] state_1_4_shl;
  wire [4:0] state_1_4_pad;
  wire [2:0] state__1_shl;
  wire [4:0] state__1_pad;
  wire [3:0] state_1_1_shl;
  wire [4:0] state_1_1_pad;
  wire [4:0] state_1_2_shl;
  wire [4:0] state_1_2_pad;
  wire [4:0] TLBroadcast_xor1;
  wire [4:0] TLBroadcast_xor6;
  wire [4:0] TLBroadcast_xor2;
  wire [4:0] TLBroadcast_xor0;
  wire [29:0] TLBroadcastTracker_sum;
  wire [29:0] TLBroadcastTracker_2_sum;
  wire [29:0] BroadcastFilter_sum;
  wire [29:0] TLBroadcastTracker_3_sum;
  wire [29:0] TLBroadcastTracker_1_sum;
  BroadcastFilter BroadcastFilter ( // @[Broadcast.scala 99:26]
    .io_request_ready(BroadcastFilter_io_request_ready),
    .io_request_valid(BroadcastFilter_io_request_valid),
    .io_response_ready(BroadcastFilter_io_response_ready),
    .io_response_valid(BroadcastFilter_io_response_valid),
    .io_covSum(BroadcastFilter_io_covSum)
  );
  TLBroadcastTracker TLBroadcastTracker ( // @[Broadcast.scala 107:15]
    .clock(TLBroadcastTracker_clock),
    .reset(TLBroadcastTracker_reset),
    .io_in_a_first(TLBroadcastTracker_io_in_a_first),
    .io_in_a_ready(TLBroadcastTracker_io_in_a_ready),
    .io_in_a_valid(TLBroadcastTracker_io_in_a_valid),
    .io_in_a_bits_opcode(TLBroadcastTracker_io_in_a_bits_opcode),
    .io_in_a_bits_size(TLBroadcastTracker_io_in_a_bits_size),
    .io_in_a_bits_source(TLBroadcastTracker_io_in_a_bits_source),
    .io_in_a_bits_address(TLBroadcastTracker_io_in_a_bits_address),
    .io_in_a_bits_user_amba_prot_bufferable(TLBroadcastTracker_io_in_a_bits_user_amba_prot_bufferable),
    .io_in_a_bits_user_amba_prot_modifiable(TLBroadcastTracker_io_in_a_bits_user_amba_prot_modifiable),
    .io_in_a_bits_user_amba_prot_readalloc(TLBroadcastTracker_io_in_a_bits_user_amba_prot_readalloc),
    .io_in_a_bits_user_amba_prot_writealloc(TLBroadcastTracker_io_in_a_bits_user_amba_prot_writealloc),
    .io_in_a_bits_user_amba_prot_privileged(TLBroadcastTracker_io_in_a_bits_user_amba_prot_privileged),
    .io_in_a_bits_user_amba_prot_secure(TLBroadcastTracker_io_in_a_bits_user_amba_prot_secure),
    .io_in_a_bits_user_amba_prot_fetch(TLBroadcastTracker_io_in_a_bits_user_amba_prot_fetch),
    .io_in_a_bits_mask(TLBroadcastTracker_io_in_a_bits_mask),
    .io_in_a_bits_data(TLBroadcastTracker_io_in_a_bits_data),
    .io_out_a_ready(TLBroadcastTracker_io_out_a_ready),
    .io_out_a_valid(TLBroadcastTracker_io_out_a_valid),
    .io_out_a_bits_opcode(TLBroadcastTracker_io_out_a_bits_opcode),
    .io_out_a_bits_size(TLBroadcastTracker_io_out_a_bits_size),
    .io_out_a_bits_source(TLBroadcastTracker_io_out_a_bits_source),
    .io_out_a_bits_address(TLBroadcastTracker_io_out_a_bits_address),
    .io_out_a_bits_user_amba_prot_bufferable(TLBroadcastTracker_io_out_a_bits_user_amba_prot_bufferable),
    .io_out_a_bits_user_amba_prot_modifiable(TLBroadcastTracker_io_out_a_bits_user_amba_prot_modifiable),
    .io_out_a_bits_user_amba_prot_readalloc(TLBroadcastTracker_io_out_a_bits_user_amba_prot_readalloc),
    .io_out_a_bits_user_amba_prot_writealloc(TLBroadcastTracker_io_out_a_bits_user_amba_prot_writealloc),
    .io_out_a_bits_user_amba_prot_privileged(TLBroadcastTracker_io_out_a_bits_user_amba_prot_privileged),
    .io_out_a_bits_user_amba_prot_secure(TLBroadcastTracker_io_out_a_bits_user_amba_prot_secure),
    .io_out_a_bits_user_amba_prot_fetch(TLBroadcastTracker_io_out_a_bits_user_amba_prot_fetch),
    .io_out_a_bits_mask(TLBroadcastTracker_io_out_a_bits_mask),
    .io_out_a_bits_data(TLBroadcastTracker_io_out_a_bits_data),
    .io_probedack(TLBroadcastTracker_io_probedack),
    .io_d_last(TLBroadcastTracker_io_d_last),
    .io_source(TLBroadcastTracker_io_source),
    .io_line(TLBroadcastTracker_io_line),
    .io_idle(TLBroadcastTracker_io_idle),
    .io_need_d(TLBroadcastTracker_io_need_d),
    .io_covSum(TLBroadcastTracker_io_covSum)
  );
  TLBroadcastTracker_1 TLBroadcastTracker_1 ( // @[Broadcast.scala 107:15]
    .clock(TLBroadcastTracker_1_clock),
    .reset(TLBroadcastTracker_1_reset),
    .io_in_a_first(TLBroadcastTracker_1_io_in_a_first),
    .io_in_a_ready(TLBroadcastTracker_1_io_in_a_ready),
    .io_in_a_valid(TLBroadcastTracker_1_io_in_a_valid),
    .io_in_a_bits_opcode(TLBroadcastTracker_1_io_in_a_bits_opcode),
    .io_in_a_bits_size(TLBroadcastTracker_1_io_in_a_bits_size),
    .io_in_a_bits_source(TLBroadcastTracker_1_io_in_a_bits_source),
    .io_in_a_bits_address(TLBroadcastTracker_1_io_in_a_bits_address),
    .io_in_a_bits_user_amba_prot_bufferable(TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_bufferable),
    .io_in_a_bits_user_amba_prot_modifiable(TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_modifiable),
    .io_in_a_bits_user_amba_prot_readalloc(TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_readalloc),
    .io_in_a_bits_user_amba_prot_writealloc(TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_writealloc),
    .io_in_a_bits_user_amba_prot_privileged(TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_privileged),
    .io_in_a_bits_user_amba_prot_secure(TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_secure),
    .io_in_a_bits_user_amba_prot_fetch(TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_fetch),
    .io_in_a_bits_mask(TLBroadcastTracker_1_io_in_a_bits_mask),
    .io_in_a_bits_data(TLBroadcastTracker_1_io_in_a_bits_data),
    .io_out_a_ready(TLBroadcastTracker_1_io_out_a_ready),
    .io_out_a_valid(TLBroadcastTracker_1_io_out_a_valid),
    .io_out_a_bits_opcode(TLBroadcastTracker_1_io_out_a_bits_opcode),
    .io_out_a_bits_size(TLBroadcastTracker_1_io_out_a_bits_size),
    .io_out_a_bits_source(TLBroadcastTracker_1_io_out_a_bits_source),
    .io_out_a_bits_address(TLBroadcastTracker_1_io_out_a_bits_address),
    .io_out_a_bits_user_amba_prot_bufferable(TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_bufferable),
    .io_out_a_bits_user_amba_prot_modifiable(TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_modifiable),
    .io_out_a_bits_user_amba_prot_readalloc(TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_readalloc),
    .io_out_a_bits_user_amba_prot_writealloc(TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_writealloc),
    .io_out_a_bits_user_amba_prot_privileged(TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_privileged),
    .io_out_a_bits_user_amba_prot_secure(TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_secure),
    .io_out_a_bits_user_amba_prot_fetch(TLBroadcastTracker_1_io_out_a_bits_user_amba_prot_fetch),
    .io_out_a_bits_mask(TLBroadcastTracker_1_io_out_a_bits_mask),
    .io_out_a_bits_data(TLBroadcastTracker_1_io_out_a_bits_data),
    .io_probedack(TLBroadcastTracker_1_io_probedack),
    .io_d_last(TLBroadcastTracker_1_io_d_last),
    .io_source(TLBroadcastTracker_1_io_source),
    .io_line(TLBroadcastTracker_1_io_line),
    .io_idle(TLBroadcastTracker_1_io_idle),
    .io_need_d(TLBroadcastTracker_1_io_need_d),
    .io_covSum(TLBroadcastTracker_1_io_covSum)
  );
  TLBroadcastTracker_2 TLBroadcastTracker_2 ( // @[Broadcast.scala 107:15]
    .clock(TLBroadcastTracker_2_clock),
    .reset(TLBroadcastTracker_2_reset),
    .io_in_a_first(TLBroadcastTracker_2_io_in_a_first),
    .io_in_a_ready(TLBroadcastTracker_2_io_in_a_ready),
    .io_in_a_valid(TLBroadcastTracker_2_io_in_a_valid),
    .io_in_a_bits_opcode(TLBroadcastTracker_2_io_in_a_bits_opcode),
    .io_in_a_bits_size(TLBroadcastTracker_2_io_in_a_bits_size),
    .io_in_a_bits_source(TLBroadcastTracker_2_io_in_a_bits_source),
    .io_in_a_bits_address(TLBroadcastTracker_2_io_in_a_bits_address),
    .io_in_a_bits_user_amba_prot_bufferable(TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_bufferable),
    .io_in_a_bits_user_amba_prot_modifiable(TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_modifiable),
    .io_in_a_bits_user_amba_prot_readalloc(TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_readalloc),
    .io_in_a_bits_user_amba_prot_writealloc(TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_writealloc),
    .io_in_a_bits_user_amba_prot_privileged(TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_privileged),
    .io_in_a_bits_user_amba_prot_secure(TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_secure),
    .io_in_a_bits_user_amba_prot_fetch(TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_fetch),
    .io_in_a_bits_mask(TLBroadcastTracker_2_io_in_a_bits_mask),
    .io_in_a_bits_data(TLBroadcastTracker_2_io_in_a_bits_data),
    .io_out_a_ready(TLBroadcastTracker_2_io_out_a_ready),
    .io_out_a_valid(TLBroadcastTracker_2_io_out_a_valid),
    .io_out_a_bits_opcode(TLBroadcastTracker_2_io_out_a_bits_opcode),
    .io_out_a_bits_size(TLBroadcastTracker_2_io_out_a_bits_size),
    .io_out_a_bits_source(TLBroadcastTracker_2_io_out_a_bits_source),
    .io_out_a_bits_address(TLBroadcastTracker_2_io_out_a_bits_address),
    .io_out_a_bits_user_amba_prot_bufferable(TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_bufferable),
    .io_out_a_bits_user_amba_prot_modifiable(TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_modifiable),
    .io_out_a_bits_user_amba_prot_readalloc(TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_readalloc),
    .io_out_a_bits_user_amba_prot_writealloc(TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_writealloc),
    .io_out_a_bits_user_amba_prot_privileged(TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_privileged),
    .io_out_a_bits_user_amba_prot_secure(TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_secure),
    .io_out_a_bits_user_amba_prot_fetch(TLBroadcastTracker_2_io_out_a_bits_user_amba_prot_fetch),
    .io_out_a_bits_mask(TLBroadcastTracker_2_io_out_a_bits_mask),
    .io_out_a_bits_data(TLBroadcastTracker_2_io_out_a_bits_data),
    .io_probedack(TLBroadcastTracker_2_io_probedack),
    .io_d_last(TLBroadcastTracker_2_io_d_last),
    .io_source(TLBroadcastTracker_2_io_source),
    .io_line(TLBroadcastTracker_2_io_line),
    .io_idle(TLBroadcastTracker_2_io_idle),
    .io_need_d(TLBroadcastTracker_2_io_need_d),
    .io_covSum(TLBroadcastTracker_2_io_covSum)
  );
  TLBroadcastTracker_3 TLBroadcastTracker_3 ( // @[Broadcast.scala 107:15]
    .clock(TLBroadcastTracker_3_clock),
    .reset(TLBroadcastTracker_3_reset),
    .io_in_a_first(TLBroadcastTracker_3_io_in_a_first),
    .io_in_a_ready(TLBroadcastTracker_3_io_in_a_ready),
    .io_in_a_valid(TLBroadcastTracker_3_io_in_a_valid),
    .io_in_a_bits_opcode(TLBroadcastTracker_3_io_in_a_bits_opcode),
    .io_in_a_bits_size(TLBroadcastTracker_3_io_in_a_bits_size),
    .io_in_a_bits_source(TLBroadcastTracker_3_io_in_a_bits_source),
    .io_in_a_bits_address(TLBroadcastTracker_3_io_in_a_bits_address),
    .io_in_a_bits_user_amba_prot_bufferable(TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_bufferable),
    .io_in_a_bits_user_amba_prot_modifiable(TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_modifiable),
    .io_in_a_bits_user_amba_prot_readalloc(TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_readalloc),
    .io_in_a_bits_user_amba_prot_writealloc(TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_writealloc),
    .io_in_a_bits_user_amba_prot_privileged(TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_privileged),
    .io_in_a_bits_user_amba_prot_secure(TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_secure),
    .io_in_a_bits_user_amba_prot_fetch(TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_fetch),
    .io_in_a_bits_mask(TLBroadcastTracker_3_io_in_a_bits_mask),
    .io_in_a_bits_data(TLBroadcastTracker_3_io_in_a_bits_data),
    .io_out_a_ready(TLBroadcastTracker_3_io_out_a_ready),
    .io_out_a_valid(TLBroadcastTracker_3_io_out_a_valid),
    .io_out_a_bits_opcode(TLBroadcastTracker_3_io_out_a_bits_opcode),
    .io_out_a_bits_size(TLBroadcastTracker_3_io_out_a_bits_size),
    .io_out_a_bits_source(TLBroadcastTracker_3_io_out_a_bits_source),
    .io_out_a_bits_address(TLBroadcastTracker_3_io_out_a_bits_address),
    .io_out_a_bits_user_amba_prot_bufferable(TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_bufferable),
    .io_out_a_bits_user_amba_prot_modifiable(TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_modifiable),
    .io_out_a_bits_user_amba_prot_readalloc(TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_readalloc),
    .io_out_a_bits_user_amba_prot_writealloc(TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_writealloc),
    .io_out_a_bits_user_amba_prot_privileged(TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_privileged),
    .io_out_a_bits_user_amba_prot_secure(TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_secure),
    .io_out_a_bits_user_amba_prot_fetch(TLBroadcastTracker_3_io_out_a_bits_user_amba_prot_fetch),
    .io_out_a_bits_mask(TLBroadcastTracker_3_io_out_a_bits_mask),
    .io_out_a_bits_data(TLBroadcastTracker_3_io_out_a_bits_data),
    .io_probedack(TLBroadcastTracker_3_io_probedack),
    .io_d_last(TLBroadcastTracker_3_io_d_last),
    .io_source(TLBroadcastTracker_3_io_source),
    .io_line(TLBroadcastTracker_3_io_line),
    .io_idle(TLBroadcastTracker_3_io_idle),
    .io_need_d(TLBroadcastTracker_3_io_need_d),
    .io_covSum(TLBroadcastTracker_3_io_covSum)
  );
  assign auto_in_a_ready = (~first_2 | BroadcastFilter_io_request_ready) & _T_478; // @[Broadcast.scala 243:59]
  assign auto_in_d_valid = idle ? out_1_earlyValid : _sink_ACancel_earlyValid_T_2; // @[Arbiter.scala 125:29]
  assign auto_in_d_bits_opcode = muxStateEarly__1 ? out_1_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  assign auto_in_d_bits_size = muxStateEarly__1 ? auto_out_d_bits_size : 3'h0; // @[Mux.scala 27:73]
  assign auto_in_d_bits_source = muxStateEarly__1 ? out_1_bits_source : 7'h0; // @[Mux.scala 27:73]
  assign auto_in_d_bits_denied = muxStateEarly__1 & auto_out_d_bits_denied; // @[Mux.scala 27:73]
  assign auto_in_d_bits_data = muxStateEarly__1 ? auto_out_d_bits_data : 64'h0; // @[Mux.scala 27:73]
  assign auto_in_d_bits_corrupt = muxStateEarly__1 & auto_out_d_bits_corrupt; // @[Mux.scala 27:73]
  assign auto_out_a_valid = idle_1 ? _T_286 : _sink_ACancel_earlyValid_T_17; // @[Arbiter.scala 125:29]
  assign auto_out_a_bits_opcode = _T_442 | _T_439; // @[Mux.scala 27:73]
  assign auto_out_a_bits_size = _T_424 | _T_421; // @[Mux.scala 27:73]
  assign auto_out_a_bits_source = _T_415 | _T_412; // @[Mux.scala 27:73]
  assign auto_out_a_bits_address = _T_406 | _T_403; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_bufferable = muxStateEarly_1_1 & out_4_bits_user_amba_prot_bufferable |
    muxStateEarly_1_2 & out_5_bits_user_amba_prot_bufferable | muxStateEarly_1_3 & out_6_bits_user_amba_prot_bufferable
     | muxStateEarly_1_4 & out_7_bits_user_amba_prot_bufferable; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_modifiable = muxStateEarly_1_1 & out_4_bits_user_amba_prot_modifiable |
    muxStateEarly_1_2 & out_5_bits_user_amba_prot_modifiable | muxStateEarly_1_3 & out_6_bits_user_amba_prot_modifiable
     | muxStateEarly_1_4 & out_7_bits_user_amba_prot_modifiable; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_readalloc = muxStateEarly_1_1 & out_4_bits_user_amba_prot_readalloc |
    muxStateEarly_1_2 & out_5_bits_user_amba_prot_readalloc | muxStateEarly_1_3 & out_6_bits_user_amba_prot_readalloc |
    muxStateEarly_1_4 & out_7_bits_user_amba_prot_readalloc; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_writealloc = muxStateEarly_1_1 & out_4_bits_user_amba_prot_writealloc |
    muxStateEarly_1_2 & out_5_bits_user_amba_prot_writealloc | muxStateEarly_1_3 & out_6_bits_user_amba_prot_writealloc
     | muxStateEarly_1_4 & out_7_bits_user_amba_prot_writealloc; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_privileged = muxStateEarly_1_1 & out_4_bits_user_amba_prot_privileged |
    muxStateEarly_1_2 & out_5_bits_user_amba_prot_privileged | muxStateEarly_1_3 & out_6_bits_user_amba_prot_privileged
     | muxStateEarly_1_4 & out_7_bits_user_amba_prot_privileged; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_secure = muxStateEarly_1_1 & out_4_bits_user_amba_prot_secure |
    muxStateEarly_1_2 & out_5_bits_user_amba_prot_secure | muxStateEarly_1_3 & out_6_bits_user_amba_prot_secure |
    muxStateEarly_1_4 & out_7_bits_user_amba_prot_secure; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_fetch = muxStateEarly_1_1 & out_4_bits_user_amba_prot_fetch | muxStateEarly_1_2
     & out_5_bits_user_amba_prot_fetch | muxStateEarly_1_3 & out_6_bits_user_amba_prot_fetch | muxStateEarly_1_4 &
    out_7_bits_user_amba_prot_fetch; // @[Mux.scala 27:73]
  assign auto_out_a_bits_mask = _T_334 | _T_331; // @[Mux.scala 27:73]
  assign auto_out_a_bits_data = _T_325 | _T_322; // @[Mux.scala 27:73]
  assign auto_out_d_ready = out_1_ready | _T_14; // @[Broadcast.scala 128:50]
  assign BroadcastFilter_io_request_valid = auto_in_a_valid & first_2 & _T_478; // @[Broadcast.scala 250:56]
  assign BroadcastFilter_io_response_ready = ~_T_448; // @[Broadcast.scala 259:35]
  assign TLBroadcastTracker_clock = clock;
  assign TLBroadcastTracker_reset = reset;
  assign TLBroadcastTracker_io_in_a_first = counter_2 == 3'h0; // @[Edges.scala 230:25]
  assign TLBroadcastTracker_io_in_a_valid = auto_in_a_valid & _T_475[0] & _bundleIn_0_a_ready_T_1; // @[Broadcast.scala 245:46]
  assign TLBroadcastTracker_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_in_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_io_out_a_ready = auto_out_a_ready & allowed_1_1; // @[Arbiter.scala 123:31]
  assign TLBroadcastTracker_io_probedack = _GEN_1[0] & _T_65 & _T_14; // @[Broadcast.scala 143:53]
  assign TLBroadcastTracker_io_d_last = _GEN_1[0] & _T_15 & _T_56 & last; // @[Broadcast.scala 142:67]
  assign TLBroadcastTracker_1_clock = clock;
  assign TLBroadcastTracker_1_reset = reset;
  assign TLBroadcastTracker_1_io_in_a_first = counter_2 == 3'h0; // @[Edges.scala 230:25]
  assign TLBroadcastTracker_1_io_in_a_valid = auto_in_a_valid & _T_475[1] & _bundleIn_0_a_ready_T_1; // @[Broadcast.scala 245:46]
  assign TLBroadcastTracker_1_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_in_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_1_io_out_a_ready = auto_out_a_ready & allowed_1_2; // @[Arbiter.scala 123:31]
  assign TLBroadcastTracker_1_io_probedack = _GEN_1[1] & _T_65 & _T_14; // @[Broadcast.scala 143:53]
  assign TLBroadcastTracker_1_io_d_last = _GEN_1[1] & _T_15 & _T_56 & last; // @[Broadcast.scala 142:67]
  assign TLBroadcastTracker_2_clock = clock;
  assign TLBroadcastTracker_2_reset = reset;
  assign TLBroadcastTracker_2_io_in_a_first = counter_2 == 3'h0; // @[Edges.scala 230:25]
  assign TLBroadcastTracker_2_io_in_a_valid = auto_in_a_valid & _T_475[2] & _bundleIn_0_a_ready_T_1; // @[Broadcast.scala 245:46]
  assign TLBroadcastTracker_2_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_in_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_2_io_out_a_ready = auto_out_a_ready & allowed_1_3; // @[Arbiter.scala 123:31]
  assign TLBroadcastTracker_2_io_probedack = _GEN_1[2] & _T_65 & _T_14; // @[Broadcast.scala 143:53]
  assign TLBroadcastTracker_2_io_d_last = _GEN_1[2] & _T_15 & _T_56 & last; // @[Broadcast.scala 142:67]
  assign TLBroadcastTracker_3_clock = clock;
  assign TLBroadcastTracker_3_reset = reset;
  assign TLBroadcastTracker_3_io_in_a_first = counter_2 == 3'h0; // @[Edges.scala 230:25]
  assign TLBroadcastTracker_3_io_in_a_valid = auto_in_a_valid & _T_475[3] & _bundleIn_0_a_ready_T_1; // @[Broadcast.scala 245:46]
  assign TLBroadcastTracker_3_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_in_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBroadcastTracker_3_io_out_a_ready = auto_out_a_ready & allowed_1_4; // @[Arbiter.scala 123:31]
  assign TLBroadcastTracker_3_io_probedack = _GEN_1[3] & _T_65 & _T_14; // @[Broadcast.scala 143:53]
  assign TLBroadcastTracker_3_io_d_last = _GEN_1[3] & _T_15 & _T_56 & last; // @[Broadcast.scala 142:67]
  assign TLBroadcast_covMap_read_en = 1'h1;
  assign TLBroadcast_covMap_read_addr = TLBroadcast_covState;
  assign TLBroadcast_covMap_read_data = TLBroadcast_covMap[TLBroadcast_covMap_read_addr]; // @[Coverage map for TLBroadcast]
  assign TLBroadcast_covMap_write_data = 1'h1;
  assign TLBroadcast_covMap_write_addr = TLBroadcast_covState;
  assign TLBroadcast_covMap_write_mask = 1'h1;
  assign TLBroadcast_covMap_write_en = ~metaReset;
  assign state_1_3_shl = state_1_3;
  assign state_1_3_pad = {4'h0,state_1_3_shl};
  assign state_1_4_shl = {state_1_4, 1'h0};
  assign state_1_4_pad = {3'h0,state_1_4_shl};
  assign state__1_shl = {state__1, 2'h0};
  assign state__1_pad = {2'h0,state__1_shl};
  assign state_1_1_shl = {state_1_1, 3'h0};
  assign state_1_1_pad = {1'h0,state_1_1_shl};
  assign state_1_2_shl = {state_1_2, 4'h0};
  assign state_1_2_pad = state_1_2_shl;
  assign TLBroadcast_xor1 = state_1_3_pad ^ state_1_4_pad;
  assign TLBroadcast_xor6 = state_1_1_pad ^ state_1_2_pad;
  assign TLBroadcast_xor2 = state__1_pad ^ TLBroadcast_xor6;
  assign TLBroadcast_xor0 = TLBroadcast_xor1 ^ TLBroadcast_xor2;
  assign TLBroadcastTracker_sum = TLBroadcast_covSum + TLBroadcastTracker_io_covSum;
  assign TLBroadcastTracker_2_sum = TLBroadcastTracker_sum + TLBroadcastTracker_2_io_covSum;
  assign BroadcastFilter_sum = TLBroadcastTracker_2_sum + BroadcastFilter_io_covSum;
  assign TLBroadcastTracker_3_sum = BroadcastFilter_sum + TLBroadcastTracker_3_io_covSum;
  assign TLBroadcastTracker_1_sum = TLBroadcastTracker_3_sum + TLBroadcastTracker_1_io_covSum;
  assign io_covSum = TLBroadcastTracker_1_sum;
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 3'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin
      if (earlyWinner__1) begin
        if (beats1_opdata) begin
          beatsLeft <= beats1_decode;
        end else begin
          beatsLeft <= 3'h0;
        end
      end else begin
        beatsLeft <= 3'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter <= 3'h0; // @[Edges.scala 228:27]
    end else if (_T_15) begin
      if (first) begin
        if (beats1_opdata) begin
          counter <= beats1_decode;
        end else begin
          counter <= 3'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state__1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state__1 <= earlyWinner__1;
    end
    if (first) begin // @[Reg.scala 17:18]
      r <= _T_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft_1 <= 3'h0; // @[Arbiter.scala 87:30]
    end else if (latch_1) begin
      beatsLeft_1 <= initBeats_1;
    end else begin
      beatsLeft_1 <= _beatsLeft_T_10;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin
      state_1_1 <= earlyWinner_1_1;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1_2 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin
      state_1_2 <= earlyWinner_1_2;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1_3 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin
      state_1_3 <= earlyWinner_1_3;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1_4 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle_1) begin
      state_1_4 <= earlyWinner_1_4;
    end
    if (reset) begin // @[Broadcast.scala 215:31]
      REG <= 1'h0; // @[Broadcast.scala 215:31]
    end else begin
      REG <= _GEN_7[0];
    end
    if (reset) begin // @[Edges.scala 228:27]
      counter_2 <= 3'h0; // @[Edges.scala 228:27]
    end else if (_T_452) begin
      if (first_2) begin
        if (beats1_opdata_2) begin
          counter_2 <= beats1_decode_2;
        end else begin
          counter_2 <= 3'h0;
        end
      end else begin
        counter_2 <= counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_d_valid | _T_35 | auto_out_d_bits_opcode == 3'h0) & ~reset) begin
          $fatal; // @[Broadcast.scala 125:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_out_d_valid | _T_35 | auto_out_d_bits_opcode == 3'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Broadcast.scala:125 assert (!out.d.valid || !d_drop || out.d.bits.opcode === TLMessages.AccessAck)\n"
            ); // @[Broadcast.scala 125:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~out_1_earlyValid | (|_GEN_1 | out_1_bits_opcode == 3'h6)) & _T_32) begin
          $fatal; // @[Broadcast.scala 137:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_32 & ~(~out_1_earlyValid | (|_GEN_1 | out_1_bits_opcode == 3'h6))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Broadcast.scala:137 assert (!d_normal.valid || (d_trackerOH.orR() || d_normal.bits.opcode === TLMessages.ReleaseAck))\n"
            ); // @[Broadcast.scala 137:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & _T_32) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_46 | earlyWinner__1) & _T_32) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_32 & ~(_T_46 | earlyWinner__1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_46 | out_1_earlyValid) & _T_32) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_32 & ~(_T_46 | out_1_earlyValid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~((~earlyWinner_1_1 | ~earlyWinner_1_2) & (~prefixOR_3 | ~earlyWinner_1_3) & (~prefixOR_4 | ~earlyWinner_1_4
          )) & _T_32) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_32 & ~((~earlyWinner_1_1 | ~earlyWinner_1_2) & (~prefixOR_3 | ~earlyWinner_1_3) & (~prefixOR_4 | ~
          earlyWinner_1_4))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(out_4_earlyValid | out_5_earlyValid | out_6_earlyValid | out_7_earlyValid) | (prefixOR_4 |
          earlyWinner_1_4)) & _T_32) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_32 & ~(~(out_4_earlyValid | out_5_earlyValid | out_6_earlyValid | out_7_earlyValid) | (prefixOR_4 |
          earlyWinner_1_4))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_287 | _T_286) & _T_32) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_32 & ~(_T_287 | _T_286)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    TLBroadcast_covState <= TLBroadcast_xor0;
    if (TLBroadcast_covMap_write_en & TLBroadcast_covMap_write_mask) begin
      TLBroadcast_covMap[TLBroadcast_covMap_write_addr] <= TLBroadcast_covMap_write_data; // @[Coverage map for TLBroadcast]
    end
    if (!(TLBroadcast_covMap_read_data | metaReset)) begin
      TLBroadcast_covSum <= TLBroadcast_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    TLBroadcast_covMap[initvar] = 0; //_12[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  state__1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  beatsLeft_1 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  state_1_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_1_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_1_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_1_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  counter_2 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  TLBroadcast_covState = 0; //_11[4:0];
  _RAND_13 = {1{`RANDOM}};
  TLBroadcast_covSum = 0; //_13[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CoherenceManagerWrapper(
  input         auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready,
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid,
  output [2:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode,
  output [2:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size,
  output [8:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source,
  output [31:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address,
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_bufferable,
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_modifiable,
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_readalloc,
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_writealloc,
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_privileged,
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_secure,
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask,
  output [63:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data,
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready,
  input         auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid,
  input  [2:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode,
  input  [2:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size,
  input  [8:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source,
  input         auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied,
  input  [63:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data,
  input         auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt,
  output        auto_coherent_jbar_in_a_ready,
  input         auto_coherent_jbar_in_a_valid,
  input  [2:0]  auto_coherent_jbar_in_a_bits_opcode,
  input  [2:0]  auto_coherent_jbar_in_a_bits_size,
  input  [6:0]  auto_coherent_jbar_in_a_bits_source,
  input  [31:0] auto_coherent_jbar_in_a_bits_address,
  input         auto_coherent_jbar_in_a_bits_user_amba_prot_bufferable,
  input         auto_coherent_jbar_in_a_bits_user_amba_prot_modifiable,
  input         auto_coherent_jbar_in_a_bits_user_amba_prot_readalloc,
  input         auto_coherent_jbar_in_a_bits_user_amba_prot_writealloc,
  input         auto_coherent_jbar_in_a_bits_user_amba_prot_privileged,
  input         auto_coherent_jbar_in_a_bits_user_amba_prot_secure,
  input         auto_coherent_jbar_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_coherent_jbar_in_a_bits_mask,
  input  [63:0] auto_coherent_jbar_in_a_bits_data,
  input         auto_coherent_jbar_in_d_ready,
  output        auto_coherent_jbar_in_d_valid,
  output [2:0]  auto_coherent_jbar_in_d_bits_opcode,
  output [2:0]  auto_coherent_jbar_in_d_bits_size,
  output [6:0]  auto_coherent_jbar_in_d_bits_source,
  output        auto_coherent_jbar_in_d_bits_denied,
  output [63:0] auto_coherent_jbar_in_d_bits_data,
  output        auto_coherent_jbar_in_d_bits_corrupt,
  input         auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock,
  input         auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset,
  input         auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock,
  input         auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset,
  output        auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock,
  output        auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_clock;
  wire  subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_reset;
  wire  subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_clock;
  wire  subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_reset;
  wire  subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_clock;
  wire  subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_reset;
  wire  subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_clock;
  wire  subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_reset;
  wire  clockGroup_auto_in_member_subsystem_l2_0_clock;
  wire  clockGroup_auto_in_member_subsystem_l2_0_reset;
  wire  clockGroup_auto_out_clock;
  wire  clockGroup_auto_out_reset;
  wire  fixedClockNode_auto_in_clock;
  wire  fixedClockNode_auto_in_reset;
  wire  fixedClockNode_auto_out_clock;
  wire  fixedClockNode_auto_out_reset;
  wire  broadcast_1_clock; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_reset; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_a_ready; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_a_valid; // @[BankedL2Params.scala 81:24]
  wire [2:0] broadcast_1_auto_in_a_bits_opcode; // @[BankedL2Params.scala 81:24]
  wire [2:0] broadcast_1_auto_in_a_bits_size; // @[BankedL2Params.scala 81:24]
  wire [6:0] broadcast_1_auto_in_a_bits_source; // @[BankedL2Params.scala 81:24]
  wire [31:0] broadcast_1_auto_in_a_bits_address; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_a_bits_user_amba_prot_bufferable; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_a_bits_user_amba_prot_modifiable; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_a_bits_user_amba_prot_readalloc; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_a_bits_user_amba_prot_writealloc; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_a_bits_user_amba_prot_privileged; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_a_bits_user_amba_prot_secure; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_a_bits_user_amba_prot_fetch; // @[BankedL2Params.scala 81:24]
  wire [7:0] broadcast_1_auto_in_a_bits_mask; // @[BankedL2Params.scala 81:24]
  wire [63:0] broadcast_1_auto_in_a_bits_data; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_d_ready; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_d_valid; // @[BankedL2Params.scala 81:24]
  wire [2:0] broadcast_1_auto_in_d_bits_opcode; // @[BankedL2Params.scala 81:24]
  wire [2:0] broadcast_1_auto_in_d_bits_size; // @[BankedL2Params.scala 81:24]
  wire [6:0] broadcast_1_auto_in_d_bits_source; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_d_bits_denied; // @[BankedL2Params.scala 81:24]
  wire [63:0] broadcast_1_auto_in_d_bits_data; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_in_d_bits_corrupt; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_a_ready; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_a_valid; // @[BankedL2Params.scala 81:24]
  wire [2:0] broadcast_1_auto_out_a_bits_opcode; // @[BankedL2Params.scala 81:24]
  wire [2:0] broadcast_1_auto_out_a_bits_size; // @[BankedL2Params.scala 81:24]
  wire [8:0] broadcast_1_auto_out_a_bits_source; // @[BankedL2Params.scala 81:24]
  wire [31:0] broadcast_1_auto_out_a_bits_address; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_a_bits_user_amba_prot_bufferable; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_a_bits_user_amba_prot_modifiable; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_a_bits_user_amba_prot_readalloc; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_a_bits_user_amba_prot_writealloc; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_a_bits_user_amba_prot_privileged; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_a_bits_user_amba_prot_secure; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_a_bits_user_amba_prot_fetch; // @[BankedL2Params.scala 81:24]
  wire [7:0] broadcast_1_auto_out_a_bits_mask; // @[BankedL2Params.scala 81:24]
  wire [63:0] broadcast_1_auto_out_a_bits_data; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_d_ready; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_d_valid; // @[BankedL2Params.scala 81:24]
  wire [2:0] broadcast_1_auto_out_d_bits_opcode; // @[BankedL2Params.scala 81:24]
  wire [2:0] broadcast_1_auto_out_d_bits_size; // @[BankedL2Params.scala 81:24]
  wire [8:0] broadcast_1_auto_out_d_bits_source; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_d_bits_denied; // @[BankedL2Params.scala 81:24]
  wire [63:0] broadcast_1_auto_out_d_bits_data; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_auto_out_d_bits_corrupt; // @[BankedL2Params.scala 81:24]
  wire [29:0] broadcast_1_io_covSum; // @[BankedL2Params.scala 81:24]
  wire  broadcast_1_metaReset; // @[BankedL2Params.scala 81:24]
  wire  coherent_jbar_auto_in_a_ready;
  wire  coherent_jbar_auto_in_a_valid;
  wire [2:0] coherent_jbar_auto_in_a_bits_opcode;
  wire [2:0] coherent_jbar_auto_in_a_bits_size;
  wire [6:0] coherent_jbar_auto_in_a_bits_source;
  wire [31:0] coherent_jbar_auto_in_a_bits_address;
  wire  coherent_jbar_auto_in_a_bits_user_amba_prot_bufferable;
  wire  coherent_jbar_auto_in_a_bits_user_amba_prot_modifiable;
  wire  coherent_jbar_auto_in_a_bits_user_amba_prot_readalloc;
  wire  coherent_jbar_auto_in_a_bits_user_amba_prot_writealloc;
  wire  coherent_jbar_auto_in_a_bits_user_amba_prot_privileged;
  wire  coherent_jbar_auto_in_a_bits_user_amba_prot_secure;
  wire  coherent_jbar_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] coherent_jbar_auto_in_a_bits_mask;
  wire [63:0] coherent_jbar_auto_in_a_bits_data;
  wire  coherent_jbar_auto_in_d_ready;
  wire  coherent_jbar_auto_in_d_valid;
  wire [2:0] coherent_jbar_auto_in_d_bits_opcode;
  wire [2:0] coherent_jbar_auto_in_d_bits_size;
  wire [6:0] coherent_jbar_auto_in_d_bits_source;
  wire  coherent_jbar_auto_in_d_bits_denied;
  wire [63:0] coherent_jbar_auto_in_d_bits_data;
  wire  coherent_jbar_auto_in_d_bits_corrupt;
  wire  coherent_jbar_auto_out_a_ready;
  wire  coherent_jbar_auto_out_a_valid;
  wire [2:0] coherent_jbar_auto_out_a_bits_opcode;
  wire [2:0] coherent_jbar_auto_out_a_bits_size;
  wire [6:0] coherent_jbar_auto_out_a_bits_source;
  wire [31:0] coherent_jbar_auto_out_a_bits_address;
  wire  coherent_jbar_auto_out_a_bits_user_amba_prot_bufferable;
  wire  coherent_jbar_auto_out_a_bits_user_amba_prot_modifiable;
  wire  coherent_jbar_auto_out_a_bits_user_amba_prot_readalloc;
  wire  coherent_jbar_auto_out_a_bits_user_amba_prot_writealloc;
  wire  coherent_jbar_auto_out_a_bits_user_amba_prot_privileged;
  wire  coherent_jbar_auto_out_a_bits_user_amba_prot_secure;
  wire  coherent_jbar_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] coherent_jbar_auto_out_a_bits_mask;
  wire [63:0] coherent_jbar_auto_out_a_bits_data;
  wire  coherent_jbar_auto_out_d_ready;
  wire  coherent_jbar_auto_out_d_valid;
  wire [2:0] coherent_jbar_auto_out_d_bits_opcode;
  wire [2:0] coherent_jbar_auto_out_d_bits_size;
  wire [6:0] coherent_jbar_auto_out_d_bits_source;
  wire  coherent_jbar_auto_out_d_bits_denied;
  wire [63:0] coherent_jbar_auto_out_d_bits_data;
  wire  coherent_jbar_auto_out_d_bits_corrupt;
  wire  binder_auto_in_a_ready; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_a_valid; // @[BankBinder.scala 67:28]
  wire [2:0] binder_auto_in_a_bits_opcode; // @[BankBinder.scala 67:28]
  wire [2:0] binder_auto_in_a_bits_size; // @[BankBinder.scala 67:28]
  wire [8:0] binder_auto_in_a_bits_source; // @[BankBinder.scala 67:28]
  wire [31:0] binder_auto_in_a_bits_address; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_a_bits_user_amba_prot_bufferable; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_a_bits_user_amba_prot_modifiable; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_a_bits_user_amba_prot_readalloc; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_a_bits_user_amba_prot_writealloc; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_a_bits_user_amba_prot_privileged; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_a_bits_user_amba_prot_secure; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_a_bits_user_amba_prot_fetch; // @[BankBinder.scala 67:28]
  wire [7:0] binder_auto_in_a_bits_mask; // @[BankBinder.scala 67:28]
  wire [63:0] binder_auto_in_a_bits_data; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_d_ready; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_d_valid; // @[BankBinder.scala 67:28]
  wire [2:0] binder_auto_in_d_bits_opcode; // @[BankBinder.scala 67:28]
  wire [2:0] binder_auto_in_d_bits_size; // @[BankBinder.scala 67:28]
  wire [8:0] binder_auto_in_d_bits_source; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_d_bits_denied; // @[BankBinder.scala 67:28]
  wire [63:0] binder_auto_in_d_bits_data; // @[BankBinder.scala 67:28]
  wire  binder_auto_in_d_bits_corrupt; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_a_ready; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_a_valid; // @[BankBinder.scala 67:28]
  wire [2:0] binder_auto_out_a_bits_opcode; // @[BankBinder.scala 67:28]
  wire [2:0] binder_auto_out_a_bits_size; // @[BankBinder.scala 67:28]
  wire [8:0] binder_auto_out_a_bits_source; // @[BankBinder.scala 67:28]
  wire [31:0] binder_auto_out_a_bits_address; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_a_bits_user_amba_prot_bufferable; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_a_bits_user_amba_prot_modifiable; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_a_bits_user_amba_prot_readalloc; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_a_bits_user_amba_prot_writealloc; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_a_bits_user_amba_prot_privileged; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_a_bits_user_amba_prot_secure; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_a_bits_user_amba_prot_fetch; // @[BankBinder.scala 67:28]
  wire [7:0] binder_auto_out_a_bits_mask; // @[BankBinder.scala 67:28]
  wire [63:0] binder_auto_out_a_bits_data; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_d_ready; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_d_valid; // @[BankBinder.scala 67:28]
  wire [2:0] binder_auto_out_d_bits_opcode; // @[BankBinder.scala 67:28]
  wire [2:0] binder_auto_out_d_bits_size; // @[BankBinder.scala 67:28]
  wire [8:0] binder_auto_out_d_bits_source; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_d_bits_denied; // @[BankBinder.scala 67:28]
  wire [63:0] binder_auto_out_d_bits_data; // @[BankBinder.scala 67:28]
  wire  binder_auto_out_d_bits_corrupt; // @[BankBinder.scala 67:28]
  wire [29:0] binder_io_covSum; // @[BankBinder.scala 67:28]
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_ready;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_size;
  wire [8:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_source;
  wire [31:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_address;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_bufferable;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_modifiable;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_readalloc;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_writealloc;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_privileged;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_secure;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_data;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_ready;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_size;
  wire [8:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_source;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_data;
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_ready;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_size;
  wire [8:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_source;
  wire [31:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_address;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_bufferable;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_modifiable;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_readalloc;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_writealloc;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_privileged;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_secure;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_data;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_ready;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_size;
  wire [8:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_source;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_data;
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_ready;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_size;
  wire [8:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_source;
  wire [31:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_address;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_bufferable;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_modifiable;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_readalloc;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_writealloc;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_privileged;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_secure;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_data;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_ready;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_size;
  wire [8:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_source;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_data;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_corrupt;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_ready;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_valid;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_size;
  wire [8:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_source;
  wire [31:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_address;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_bufferable;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_modifiable;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_readalloc;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_writealloc;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_privileged;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_secure;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_mask;
  wire [63:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_data;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_ready;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_valid;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_opcode;
  wire [2:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_size;
  wire [8:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_source;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_denied;
  wire [63:0] coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_data;
  wire  coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_corrupt;
  wire [29:0] CoherenceManagerWrapper_covSum;
  wire [29:0] broadcast_1_sum;
  wire [29:0] binder_sum;
  TLBroadcast broadcast_1 ( // @[BankedL2Params.scala 81:24]
    .clock(broadcast_1_clock),
    .reset(broadcast_1_reset),
    .auto_in_a_ready(broadcast_1_auto_in_a_ready),
    .auto_in_a_valid(broadcast_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(broadcast_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(broadcast_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(broadcast_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(broadcast_1_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(broadcast_1_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(broadcast_1_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(broadcast_1_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(broadcast_1_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(broadcast_1_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(broadcast_1_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(broadcast_1_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(broadcast_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(broadcast_1_auto_in_a_bits_data),
    .auto_in_d_ready(broadcast_1_auto_in_d_ready),
    .auto_in_d_valid(broadcast_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(broadcast_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(broadcast_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(broadcast_1_auto_in_d_bits_source),
    .auto_in_d_bits_denied(broadcast_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(broadcast_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(broadcast_1_auto_in_d_bits_corrupt),
    .auto_out_a_ready(broadcast_1_auto_out_a_ready),
    .auto_out_a_valid(broadcast_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(broadcast_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(broadcast_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(broadcast_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(broadcast_1_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(broadcast_1_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(broadcast_1_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(broadcast_1_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(broadcast_1_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(broadcast_1_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(broadcast_1_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(broadcast_1_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(broadcast_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(broadcast_1_auto_out_a_bits_data),
    .auto_out_d_ready(broadcast_1_auto_out_d_ready),
    .auto_out_d_valid(broadcast_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(broadcast_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(broadcast_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(broadcast_1_auto_out_d_bits_source),
    .auto_out_d_bits_denied(broadcast_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(broadcast_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(broadcast_1_auto_out_d_bits_corrupt),
    .io_covSum(broadcast_1_io_covSum),
    .metaReset(broadcast_1_metaReset)
  );
  ProbePicker binder ( // @[BankBinder.scala 67:28]
    .auto_in_a_ready(binder_auto_in_a_ready),
    .auto_in_a_valid(binder_auto_in_a_valid),
    .auto_in_a_bits_opcode(binder_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(binder_auto_in_a_bits_size),
    .auto_in_a_bits_source(binder_auto_in_a_bits_source),
    .auto_in_a_bits_address(binder_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(binder_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(binder_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(binder_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(binder_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(binder_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(binder_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(binder_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(binder_auto_in_a_bits_mask),
    .auto_in_a_bits_data(binder_auto_in_a_bits_data),
    .auto_in_d_ready(binder_auto_in_d_ready),
    .auto_in_d_valid(binder_auto_in_d_valid),
    .auto_in_d_bits_opcode(binder_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(binder_auto_in_d_bits_size),
    .auto_in_d_bits_source(binder_auto_in_d_bits_source),
    .auto_in_d_bits_denied(binder_auto_in_d_bits_denied),
    .auto_in_d_bits_data(binder_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(binder_auto_in_d_bits_corrupt),
    .auto_out_a_ready(binder_auto_out_a_ready),
    .auto_out_a_valid(binder_auto_out_a_valid),
    .auto_out_a_bits_opcode(binder_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(binder_auto_out_a_bits_size),
    .auto_out_a_bits_source(binder_auto_out_a_bits_source),
    .auto_out_a_bits_address(binder_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(binder_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(binder_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(binder_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(binder_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(binder_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(binder_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(binder_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(binder_auto_out_a_bits_mask),
    .auto_out_a_bits_data(binder_auto_out_a_bits_data),
    .auto_out_d_ready(binder_auto_out_d_ready),
    .auto_out_d_valid(binder_auto_out_d_valid),
    .auto_out_d_bits_opcode(binder_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(binder_auto_out_d_bits_size),
    .auto_out_d_bits_source(binder_auto_out_d_bits_source),
    .auto_out_d_bits_denied(binder_auto_out_d_bits_denied),
    .auto_out_d_bits_data(binder_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(binder_auto_out_d_bits_corrupt),
    .io_covSum(binder_io_covSum)
  );
  assign subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_clock =
    subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_reset =
    subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_clock =
    subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_reset =
    subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_clock = clockGroup_auto_in_member_subsystem_l2_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockGroup_auto_out_reset = clockGroup_auto_in_member_subsystem_l2_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fixedClockNode_auto_out_clock = fixedClockNode_auto_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign fixedClockNode_auto_out_reset = fixedClockNode_auto_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_ready = coherent_jbar_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coherent_jbar_auto_in_d_valid = coherent_jbar_auto_out_d_valid; // @[ReadyValidCancel.scala 21:38]
  assign coherent_jbar_auto_in_d_bits_opcode = coherent_jbar_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coherent_jbar_auto_in_d_bits_size = coherent_jbar_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coherent_jbar_auto_in_d_bits_source = coherent_jbar_auto_out_d_bits_source; // @[Xbar.scala 228:69]
  assign coherent_jbar_auto_in_d_bits_denied = coherent_jbar_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coherent_jbar_auto_in_d_bits_data = coherent_jbar_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coherent_jbar_auto_in_d_bits_corrupt = coherent_jbar_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coherent_jbar_auto_out_a_valid = coherent_jbar_auto_in_a_valid; // @[ReadyValidCancel.scala 21:38]
  assign coherent_jbar_auto_out_a_bits_opcode = coherent_jbar_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_size = coherent_jbar_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_source = coherent_jbar_auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign coherent_jbar_auto_out_a_bits_address = coherent_jbar_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_user_amba_prot_bufferable =
    coherent_jbar_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_user_amba_prot_modifiable =
    coherent_jbar_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_user_amba_prot_readalloc = coherent_jbar_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_user_amba_prot_writealloc =
    coherent_jbar_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_user_amba_prot_privileged =
    coherent_jbar_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_user_amba_prot_secure = coherent_jbar_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_user_amba_prot_fetch = coherent_jbar_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_mask = coherent_jbar_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_bits_data = coherent_jbar_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_d_ready = coherent_jbar_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_ready =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_valid =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_opcode =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_size =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_source =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_denied =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_data =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_corrupt =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_valid =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_size =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_source =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_address =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_bufferable =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_modifiable =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_readalloc =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_writealloc =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_privileged =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_secure =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_fetch =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_mask =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_data =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_ready =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_ready =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_ready; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_valid =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_valid; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_opcode =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_size =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_source =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_denied =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_denied; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_data =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_corrupt =
    coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_valid =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_size =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_source =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_address =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_bufferable =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_modifiable =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_readalloc =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_writealloc =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_privileged =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_secure =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_fetch =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_mask =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_data =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_ready =
    coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_valid =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_valid; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_opcode =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_size =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_source =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_address =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_bufferable =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_modifiable =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_readalloc =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_writealloc =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_privileged =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_secure =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_secure; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_user_amba_prot_fetch =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_mask =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_a_bits_data =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_in_d_ready =
    coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_ready; // @[LazyModule.scala 309:16]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_a_ready =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_valid =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_opcode =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_size =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_source =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_denied =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_data =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_widget_auto_out_d_bits_corrupt =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_bufferable =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_modifiable =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_readalloc =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_writealloc =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_privileged =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_secure =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_fetch =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_coherent_jbar_in_a_ready = coherent_jbar_auto_in_a_ready; // @[LazyModule.scala 309:16]
  assign auto_coherent_jbar_in_d_valid = coherent_jbar_auto_in_d_valid; // @[LazyModule.scala 309:16]
  assign auto_coherent_jbar_in_d_bits_opcode = coherent_jbar_auto_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign auto_coherent_jbar_in_d_bits_size = coherent_jbar_auto_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_coherent_jbar_in_d_bits_source = coherent_jbar_auto_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign auto_coherent_jbar_in_d_bits_denied = coherent_jbar_auto_in_d_bits_denied; // @[LazyModule.scala 309:16]
  assign auto_coherent_jbar_in_d_bits_data = coherent_jbar_auto_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign auto_coherent_jbar_in_d_bits_corrupt = coherent_jbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock =
    subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_clock; // @[LazyModule.scala 311:12]
  assign auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset =
    subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_reset; // @[LazyModule.scala 311:12]
  assign subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_clock =
    auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock; // @[LazyModule.scala 309:16]
  assign subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_reset =
    auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset; // @[LazyModule.scala 309:16]
  assign subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_clock =
    auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock; // @[LazyModule.scala 309:16]
  assign subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_reset =
    auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset; // @[LazyModule.scala 309:16]
  assign clockGroup_auto_in_member_subsystem_l2_0_clock =
    subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_clock; // @[LazyModule.scala 298:16]
  assign clockGroup_auto_in_member_subsystem_l2_0_reset =
    subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_reset; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[LazyModule.scala 298:16]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[LazyModule.scala 298:16]
  assign broadcast_1_clock = fixedClockNode_auto_out_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign broadcast_1_reset = fixedClockNode_auto_out_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_valid = coherent_jbar_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_opcode = coherent_jbar_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_size = coherent_jbar_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_source = coherent_jbar_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_address = coherent_jbar_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_user_amba_prot_bufferable = coherent_jbar_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_user_amba_prot_modifiable = coherent_jbar_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_user_amba_prot_readalloc = coherent_jbar_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_user_amba_prot_writealloc = coherent_jbar_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_user_amba_prot_privileged = coherent_jbar_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_user_amba_prot_secure = coherent_jbar_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_user_amba_prot_fetch = coherent_jbar_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_mask = coherent_jbar_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_a_bits_data = coherent_jbar_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_in_d_ready = coherent_jbar_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign broadcast_1_auto_out_a_ready = binder_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign broadcast_1_auto_out_d_valid = binder_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign broadcast_1_auto_out_d_bits_opcode = binder_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign broadcast_1_auto_out_d_bits_size = binder_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign broadcast_1_auto_out_d_bits_source = binder_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign broadcast_1_auto_out_d_bits_denied = binder_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign broadcast_1_auto_out_d_bits_data = binder_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign broadcast_1_auto_out_d_bits_corrupt = binder_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign coherent_jbar_auto_in_a_valid = auto_coherent_jbar_in_a_valid; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_opcode = auto_coherent_jbar_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_size = auto_coherent_jbar_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_source = auto_coherent_jbar_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_address = auto_coherent_jbar_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_user_amba_prot_bufferable = auto_coherent_jbar_in_a_bits_user_amba_prot_bufferable
    ; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_user_amba_prot_modifiable = auto_coherent_jbar_in_a_bits_user_amba_prot_modifiable
    ; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_user_amba_prot_readalloc = auto_coherent_jbar_in_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_user_amba_prot_writealloc = auto_coherent_jbar_in_a_bits_user_amba_prot_writealloc
    ; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_user_amba_prot_privileged = auto_coherent_jbar_in_a_bits_user_amba_prot_privileged
    ; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_user_amba_prot_secure = auto_coherent_jbar_in_a_bits_user_amba_prot_secure; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_user_amba_prot_fetch = auto_coherent_jbar_in_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_mask = auto_coherent_jbar_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_a_bits_data = auto_coherent_jbar_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_in_d_ready = auto_coherent_jbar_in_d_ready; // @[LazyModule.scala 309:16]
  assign coherent_jbar_auto_out_a_ready = broadcast_1_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign coherent_jbar_auto_out_d_valid = broadcast_1_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign coherent_jbar_auto_out_d_bits_opcode = broadcast_1_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign coherent_jbar_auto_out_d_bits_size = broadcast_1_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign coherent_jbar_auto_out_d_bits_source = broadcast_1_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign coherent_jbar_auto_out_d_bits_denied = broadcast_1_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign coherent_jbar_auto_out_d_bits_data = broadcast_1_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign coherent_jbar_auto_out_d_bits_corrupt = broadcast_1_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign binder_auto_in_a_valid = broadcast_1_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_opcode = broadcast_1_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_size = broadcast_1_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_source = broadcast_1_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_address = broadcast_1_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_user_amba_prot_bufferable = broadcast_1_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_user_amba_prot_modifiable = broadcast_1_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_user_amba_prot_readalloc = broadcast_1_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_user_amba_prot_writealloc = broadcast_1_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_user_amba_prot_privileged = broadcast_1_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_user_amba_prot_secure = broadcast_1_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_user_amba_prot_fetch = broadcast_1_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_mask = broadcast_1_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign binder_auto_in_a_bits_data = broadcast_1_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign binder_auto_in_d_ready = broadcast_1_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign binder_auto_out_a_ready = coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_ready; // @[LazyModule.scala 298:16]
  assign binder_auto_out_d_valid = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_valid; // @[LazyModule.scala 298:16]
  assign binder_auto_out_d_bits_opcode = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign binder_auto_out_d_bits_size = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign binder_auto_out_d_bits_source = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign binder_auto_out_d_bits_denied = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign binder_auto_out_d_bits_data = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign binder_auto_out_d_bits_corrupt = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_valid = binder_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_opcode = binder_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_size = binder_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_source = binder_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_address = binder_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_bufferable =
    binder_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_modifiable =
    binder_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_readalloc =
    binder_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_writealloc =
    binder_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_privileged =
    binder_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_secure =
    binder_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_user_amba_prot_fetch =
    binder_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_mask = binder_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_data = binder_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_ready = binder_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_ready =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_valid =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_opcode =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_size =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_source =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_denied =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_data =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_corrupt =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign CoherenceManagerWrapper_covSum = 30'h0;
  assign broadcast_1_sum = CoherenceManagerWrapper_covSum + broadcast_1_io_covSum;
  assign binder_sum = broadcast_1_sum + binder_io_covSum;
  assign io_covSum = binder_sum;
  assign broadcast_1_metaReset = metaReset;
endmodule
module IntXbar_1(
  input         auto_int_in_3_0,
  input         auto_int_in_2_0,
  input         auto_int_in_1_0,
  input         auto_int_in_1_1,
  output        auto_int_out_1,
  output        auto_int_out_2,
  output        auto_int_out_3,
  output        auto_int_out_4,
  output [29:0] io_covSum
);
  wire [29:0] IntXbar_1_covSum;
  assign auto_int_out_1 = auto_int_in_1_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_int_out_2 = auto_int_in_1_1; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_int_out_3 = auto_int_in_2_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_int_out_4 = auto_int_in_3_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign IntXbar_1_covSum = 30'h0;
  assign io_covSum = IntXbar_1_covSum;
endmodule
module Queue_24(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [5:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input         io_enq_bits_user_amba_prot_bufferable,
  input         io_enq_bits_user_amba_prot_modifiable,
  input         io_enq_bits_user_amba_prot_readalloc,
  input         io_enq_bits_user_amba_prot_writealloc,
  input         io_enq_bits_user_amba_prot_privileged,
  input         io_enq_bits_user_amba_prot_secure,
  input         io_enq_bits_user_amba_prot_fetch,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [5:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output        io_deq_bits_user_amba_prot_bufferable,
  output        io_deq_bits_user_amba_prot_modifiable,
  output        io_deq_bits_user_amba_prot_readalloc,
  output        io_deq_bits_user_amba_prot_writealloc,
  output        io_deq_bits_user_amba_prot_privileged,
  output        io_deq_bits_user_amba_prot_secure,
  output        io_deq_bits_user_amba_prot_fetch,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_param_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [5:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_bufferable [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_bufferable_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_modifiable [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_modifiable_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_readalloc [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_readalloc_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_writealloc [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_writealloc_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_privileged [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_privileged_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_secure [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_secure_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_user_amba_prot_fetch [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_user_amba_prot_fetch_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_24_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_en = 1'h1;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_bufferable_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_bufferable_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_bufferable_io_deq_bits_MPORT_data =
    ram_user_amba_prot_bufferable[ram_user_amba_prot_bufferable_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_bufferable_MPORT_data = io_enq_bits_user_amba_prot_bufferable;
  assign ram_user_amba_prot_bufferable_MPORT_addr = value;
  assign ram_user_amba_prot_bufferable_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_bufferable_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_modifiable_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_modifiable_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_modifiable_io_deq_bits_MPORT_data =
    ram_user_amba_prot_modifiable[ram_user_amba_prot_modifiable_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_modifiable_MPORT_data = io_enq_bits_user_amba_prot_modifiable;
  assign ram_user_amba_prot_modifiable_MPORT_addr = value;
  assign ram_user_amba_prot_modifiable_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_modifiable_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_readalloc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_readalloc_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_readalloc_io_deq_bits_MPORT_data =
    ram_user_amba_prot_readalloc[ram_user_amba_prot_readalloc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_readalloc_MPORT_data = io_enq_bits_user_amba_prot_readalloc;
  assign ram_user_amba_prot_readalloc_MPORT_addr = value;
  assign ram_user_amba_prot_readalloc_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_readalloc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_writealloc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_writealloc_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_writealloc_io_deq_bits_MPORT_data =
    ram_user_amba_prot_writealloc[ram_user_amba_prot_writealloc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_writealloc_MPORT_data = io_enq_bits_user_amba_prot_writealloc;
  assign ram_user_amba_prot_writealloc_MPORT_addr = value;
  assign ram_user_amba_prot_writealloc_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_writealloc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_privileged_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_privileged_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_privileged_io_deq_bits_MPORT_data =
    ram_user_amba_prot_privileged[ram_user_amba_prot_privileged_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_privileged_MPORT_data = io_enq_bits_user_amba_prot_privileged;
  assign ram_user_amba_prot_privileged_MPORT_addr = value;
  assign ram_user_amba_prot_privileged_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_privileged_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_secure_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_secure_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_secure_io_deq_bits_MPORT_data =
    ram_user_amba_prot_secure[ram_user_amba_prot_secure_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_secure_MPORT_data = io_enq_bits_user_amba_prot_secure;
  assign ram_user_amba_prot_secure_MPORT_addr = value;
  assign ram_user_amba_prot_secure_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_secure_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_user_amba_prot_fetch_io_deq_bits_MPORT_en = 1'h1;
  assign ram_user_amba_prot_fetch_io_deq_bits_MPORT_addr = value_1;
  assign ram_user_amba_prot_fetch_io_deq_bits_MPORT_data =
    ram_user_amba_prot_fetch[ram_user_amba_prot_fetch_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_user_amba_prot_fetch_MPORT_data = io_enq_bits_user_amba_prot_fetch;
  assign ram_user_amba_prot_fetch_MPORT_addr = value;
  assign ram_user_amba_prot_fetch_MPORT_mask = 1'h1;
  assign ram_user_amba_prot_fetch_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_bufferable = ram_user_amba_prot_bufferable_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_modifiable = ram_user_amba_prot_modifiable_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_readalloc = ram_user_amba_prot_readalloc_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_writealloc = ram_user_amba_prot_writealloc_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_privileged = ram_user_amba_prot_privileged_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_secure = ram_user_amba_prot_secure_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_user_amba_prot_fetch = ram_user_amba_prot_fetch_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_24_covSum = 30'h0;
  assign io_covSum = Queue_24_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_bufferable_MPORT_en & ram_user_amba_prot_bufferable_MPORT_mask) begin
      ram_user_amba_prot_bufferable[ram_user_amba_prot_bufferable_MPORT_addr] <=
        ram_user_amba_prot_bufferable_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_modifiable_MPORT_en & ram_user_amba_prot_modifiable_MPORT_mask) begin
      ram_user_amba_prot_modifiable[ram_user_amba_prot_modifiable_MPORT_addr] <=
        ram_user_amba_prot_modifiable_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_readalloc_MPORT_en & ram_user_amba_prot_readalloc_MPORT_mask) begin
      ram_user_amba_prot_readalloc[ram_user_amba_prot_readalloc_MPORT_addr] <= ram_user_amba_prot_readalloc_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_writealloc_MPORT_en & ram_user_amba_prot_writealloc_MPORT_mask) begin
      ram_user_amba_prot_writealloc[ram_user_amba_prot_writealloc_MPORT_addr] <=
        ram_user_amba_prot_writealloc_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_privileged_MPORT_en & ram_user_amba_prot_privileged_MPORT_mask) begin
      ram_user_amba_prot_privileged[ram_user_amba_prot_privileged_MPORT_addr] <=
        ram_user_amba_prot_privileged_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_secure_MPORT_en & ram_user_amba_prot_secure_MPORT_mask) begin
      ram_user_amba_prot_secure[ram_user_amba_prot_secure_MPORT_addr] <= ram_user_amba_prot_secure_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_user_amba_prot_fetch_MPORT_en & ram_user_amba_prot_fetch_MPORT_mask) begin
      ram_user_amba_prot_fetch[ram_user_amba_prot_fetch_MPORT_addr] <= ram_user_amba_prot_fetch_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= value_1 + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_bufferable[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_modifiable[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_readalloc[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_writealloc[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_privileged[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_secure[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user_amba_prot_fetch[initvar] = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_12[7:0];
  _RAND_13 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_13[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  value = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  value_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  maybe_full = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_25(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [3:0]  io_enq_bits_size,
  input  [5:0]  io_enq_bits_source,
  input         io_enq_bits_denied,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_corrupt,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [3:0]  io_deq_bits_size,
  output [5:0]  io_deq_bits_source,
  output        io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_corrupt,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] ram_source [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [5:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_denied [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 259:95]
  reg  value; // @[Counter.scala 62:40]
  reg  value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_25_covSum;
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_25_covSum = 30'h0;
  assign io_covSum = Queue_25_covSum;
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      value <= value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      value_1 <= value_1 + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_5[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  value_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_8(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [2:0]  auto_in_a_bits_param,
  input  [3:0]  auto_in_a_bits_size,
  input  [5:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input         auto_in_a_bits_user_amba_prot_bufferable,
  input         auto_in_a_bits_user_amba_prot_modifiable,
  input         auto_in_a_bits_user_amba_prot_readalloc,
  input         auto_in_a_bits_user_amba_prot_writealloc,
  input         auto_in_a_bits_user_amba_prot_privileged,
  input         auto_in_a_bits_user_amba_prot_secure,
  input         auto_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [5:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [5:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output        auto_out_a_bits_user_amba_prot_bufferable,
  output        auto_out_a_bits_user_amba_prot_modifiable,
  output        auto_out_a_bits_user_amba_prot_readalloc,
  output        auto_out_a_bits_user_amba_prot_writealloc,
  output        auto_out_a_bits_user_amba_prot_privileged,
  output        auto_out_a_bits_user_amba_prot_secure,
  output        auto_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [5:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum
);
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_param; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [5:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire [31:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_bufferable; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_modifiable; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_readalloc; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_writealloc; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_privileged; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_secure; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_enq_bits_user_amba_prot_fetch; // @[Decoupled.scala 361:21]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 361:21]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [5:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [31:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_bufferable; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_modifiable; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_readalloc; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_writealloc; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_privileged; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_secure; // @[Decoupled.scala 361:21]
  wire  bundleOut_0_a_q_io_deq_bits_user_amba_prot_fetch; // @[Decoupled.scala 361:21]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [29:0] bundleOut_0_a_q_io_covSum; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [5:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [5:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 361:21]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 361:21]
  wire [29:0] bundleIn_0_d_q_io_covSum; // @[Decoupled.scala 361:21]
  wire [29:0] TLBuffer_8_covSum;
  wire [29:0] bundleOut_0_a_q_sum;
  wire [29:0] bundleIn_0_d_q_sum;
  Queue_24 bundleOut_0_a_q ( // @[Decoupled.scala 361:21]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_user_amba_prot_bufferable(bundleOut_0_a_q_io_enq_bits_user_amba_prot_bufferable),
    .io_enq_bits_user_amba_prot_modifiable(bundleOut_0_a_q_io_enq_bits_user_amba_prot_modifiable),
    .io_enq_bits_user_amba_prot_readalloc(bundleOut_0_a_q_io_enq_bits_user_amba_prot_readalloc),
    .io_enq_bits_user_amba_prot_writealloc(bundleOut_0_a_q_io_enq_bits_user_amba_prot_writealloc),
    .io_enq_bits_user_amba_prot_privileged(bundleOut_0_a_q_io_enq_bits_user_amba_prot_privileged),
    .io_enq_bits_user_amba_prot_secure(bundleOut_0_a_q_io_enq_bits_user_amba_prot_secure),
    .io_enq_bits_user_amba_prot_fetch(bundleOut_0_a_q_io_enq_bits_user_amba_prot_fetch),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_user_amba_prot_bufferable(bundleOut_0_a_q_io_deq_bits_user_amba_prot_bufferable),
    .io_deq_bits_user_amba_prot_modifiable(bundleOut_0_a_q_io_deq_bits_user_amba_prot_modifiable),
    .io_deq_bits_user_amba_prot_readalloc(bundleOut_0_a_q_io_deq_bits_user_amba_prot_readalloc),
    .io_deq_bits_user_amba_prot_writealloc(bundleOut_0_a_q_io_deq_bits_user_amba_prot_writealloc),
    .io_deq_bits_user_amba_prot_privileged(bundleOut_0_a_q_io_deq_bits_user_amba_prot_privileged),
    .io_deq_bits_user_amba_prot_secure(bundleOut_0_a_q_io_deq_bits_user_amba_prot_secure),
    .io_deq_bits_user_amba_prot_fetch(bundleOut_0_a_q_io_deq_bits_user_amba_prot_fetch),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_covSum(bundleOut_0_a_q_io_covSum)
  );
  Queue_25 bundleIn_0_d_q ( // @[Decoupled.scala 361:21]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt),
    .io_covSum(bundleIn_0_d_q_io_covSum)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 Buffer.scala 38:13]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_bufferable = bundleOut_0_a_q_io_deq_bits_user_amba_prot_bufferable; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_modifiable = bundleOut_0_a_q_io_deq_bits_user_amba_prot_modifiable; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_readalloc = bundleOut_0_a_q_io_deq_bits_user_amba_prot_readalloc; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_writealloc = bundleOut_0_a_q_io_deq_bits_user_amba_prot_writealloc; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_privileged = bundleOut_0_a_q_io_deq_bits_user_amba_prot_privileged; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_secure = bundleOut_0_a_q_io_deq_bits_user_amba_prot_secure; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_user_amba_prot_fetch = bundleOut_0_a_q_io_deq_bits_user_amba_prot_fetch; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 Buffer.scala 37:13]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 Decoupled.scala 365:17]
  assign bundleOut_0_a_q_clock = clock;
  assign bundleOut_0_a_q_reset = reset;
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_clock = clock;
  assign bundleIn_0_d_q_reset = reset;
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLBuffer_8_covSum = 30'h0;
  assign bundleOut_0_a_q_sum = TLBuffer_8_covSum + bundleOut_0_a_q_io_covSum;
  assign bundleIn_0_d_q_sum = bundleOut_0_a_q_sum + bundleIn_0_d_q_io_covSum;
  assign io_covSum = bundleIn_0_d_q_sum;
endmodule
module TLFIFOFixer_5(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [3:0]  auto_in_a_bits_size,
  input  [5:0]  auto_in_a_bits_source,
  input  [31:0] auto_in_a_bits_address,
  input         auto_in_a_bits_user_amba_prot_bufferable,
  input         auto_in_a_bits_user_amba_prot_modifiable,
  input         auto_in_a_bits_user_amba_prot_readalloc,
  input         auto_in_a_bits_user_amba_prot_writealloc,
  input         auto_in_a_bits_user_amba_prot_privileged,
  input         auto_in_a_bits_user_amba_prot_secure,
  input         auto_in_a_bits_user_amba_prot_fetch,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [3:0]  auto_in_d_bits_size,
  output [5:0]  auto_in_d_bits_source,
  output        auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output        auto_in_d_bits_corrupt,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [3:0]  auto_out_a_bits_size,
  output [5:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output        auto_out_a_bits_user_amba_prot_bufferable,
  output        auto_out_a_bits_user_amba_prot_modifiable,
  output        auto_out_a_bits_user_amba_prot_readalloc,
  output        auto_out_a_bits_user_amba_prot_writealloc,
  output        auto_out_a_bits_user_amba_prot_privileged,
  output        auto_out_a_bits_user_amba_prot_secure,
  output        auto_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [5:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_83;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_84;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] _a_id_T_1 = {1'b0,$signed(auto_in_a_bits_address)}; // @[Parameters.scala 137:49]
  wire [32:0] _a_id_T_3 = $signed(_a_id_T_1) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  a_id = $signed(_a_id_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire  a_noDomain = ~a_id; // @[FIFOFixer.scala 55:29]
  wire  stalls_a_sel = auto_in_a_bits_source[5:2] == 4'h0; // @[Parameters.scala 54:32]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25]
  reg  flight_0; // @[FIFOFixer.scala 71:27]
  reg  flight_1; // @[FIFOFixer.scala 71:27]
  reg  flight_2; // @[FIFOFixer.scala 71:27]
  reg  flight_3; // @[FIFOFixer.scala 71:27]
  reg  stalls_id; // @[Reg.scala 16:16]
  wire  stalls_0 = stalls_a_sel & a_first & (flight_0 | flight_1 | flight_2 | flight_3) & (a_noDomain | stalls_id !=
    a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_1 = auto_in_a_bits_source[5:2] == 4'h1; // @[Parameters.scala 54:32]
  reg  flight_4; // @[FIFOFixer.scala 71:27]
  reg  flight_5; // @[FIFOFixer.scala 71:27]
  reg  flight_6; // @[FIFOFixer.scala 71:27]
  reg  flight_7; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_1; // @[Reg.scala 16:16]
  wire  stalls_1 = stalls_a_sel_1 & a_first & (flight_4 | flight_5 | flight_6 | flight_7) & (a_noDomain | stalls_id_1
     != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_2 = auto_in_a_bits_source[5:2] == 4'h2; // @[Parameters.scala 54:32]
  reg  flight_8; // @[FIFOFixer.scala 71:27]
  reg  flight_9; // @[FIFOFixer.scala 71:27]
  reg  flight_10; // @[FIFOFixer.scala 71:27]
  reg  flight_11; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_2; // @[Reg.scala 16:16]
  wire  stalls_2 = stalls_a_sel_2 & a_first & (flight_8 | flight_9 | flight_10 | flight_11) & (a_noDomain | stalls_id_2
     != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_3 = auto_in_a_bits_source[5:2] == 4'h3; // @[Parameters.scala 54:32]
  reg  flight_12; // @[FIFOFixer.scala 71:27]
  reg  flight_13; // @[FIFOFixer.scala 71:27]
  reg  flight_14; // @[FIFOFixer.scala 71:27]
  reg  flight_15; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_3; // @[Reg.scala 16:16]
  wire  stalls_3 = stalls_a_sel_3 & a_first & (flight_12 | flight_13 | flight_14 | flight_15) & (a_noDomain |
    stalls_id_3 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_4 = auto_in_a_bits_source[5:2] == 4'h4; // @[Parameters.scala 54:32]
  reg  flight_16; // @[FIFOFixer.scala 71:27]
  reg  flight_17; // @[FIFOFixer.scala 71:27]
  reg  flight_18; // @[FIFOFixer.scala 71:27]
  reg  flight_19; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_4; // @[Reg.scala 16:16]
  wire  stalls_4 = stalls_a_sel_4 & a_first & (flight_16 | flight_17 | flight_18 | flight_19) & (a_noDomain |
    stalls_id_4 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_5 = auto_in_a_bits_source[5:2] == 4'h5; // @[Parameters.scala 54:32]
  reg  flight_20; // @[FIFOFixer.scala 71:27]
  reg  flight_21; // @[FIFOFixer.scala 71:27]
  reg  flight_22; // @[FIFOFixer.scala 71:27]
  reg  flight_23; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_5; // @[Reg.scala 16:16]
  wire  stalls_5 = stalls_a_sel_5 & a_first & (flight_20 | flight_21 | flight_22 | flight_23) & (a_noDomain |
    stalls_id_5 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_6 = auto_in_a_bits_source[5:2] == 4'h6; // @[Parameters.scala 54:32]
  reg  flight_24; // @[FIFOFixer.scala 71:27]
  reg  flight_25; // @[FIFOFixer.scala 71:27]
  reg  flight_26; // @[FIFOFixer.scala 71:27]
  reg  flight_27; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_6; // @[Reg.scala 16:16]
  wire  stalls_6 = stalls_a_sel_6 & a_first & (flight_24 | flight_25 | flight_26 | flight_27) & (a_noDomain |
    stalls_id_6 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_7 = auto_in_a_bits_source[5:2] == 4'h7; // @[Parameters.scala 54:32]
  reg  flight_28; // @[FIFOFixer.scala 71:27]
  reg  flight_29; // @[FIFOFixer.scala 71:27]
  reg  flight_30; // @[FIFOFixer.scala 71:27]
  reg  flight_31; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_7; // @[Reg.scala 16:16]
  wire  stalls_7 = stalls_a_sel_7 & a_first & (flight_28 | flight_29 | flight_30 | flight_31) & (a_noDomain |
    stalls_id_7 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_8 = auto_in_a_bits_source[5:2] == 4'h8; // @[Parameters.scala 54:32]
  reg  flight_32; // @[FIFOFixer.scala 71:27]
  reg  flight_33; // @[FIFOFixer.scala 71:27]
  reg  flight_34; // @[FIFOFixer.scala 71:27]
  reg  flight_35; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_8; // @[Reg.scala 16:16]
  wire  stalls_8 = stalls_a_sel_8 & a_first & (flight_32 | flight_33 | flight_34 | flight_35) & (a_noDomain |
    stalls_id_8 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_9 = auto_in_a_bits_source[5:2] == 4'h9; // @[Parameters.scala 54:32]
  reg  flight_36; // @[FIFOFixer.scala 71:27]
  reg  flight_37; // @[FIFOFixer.scala 71:27]
  reg  flight_38; // @[FIFOFixer.scala 71:27]
  reg  flight_39; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_9; // @[Reg.scala 16:16]
  wire  stalls_9 = stalls_a_sel_9 & a_first & (flight_36 | flight_37 | flight_38 | flight_39) & (a_noDomain |
    stalls_id_9 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_10 = auto_in_a_bits_source[5:2] == 4'ha; // @[Parameters.scala 54:32]
  reg  flight_40; // @[FIFOFixer.scala 71:27]
  reg  flight_41; // @[FIFOFixer.scala 71:27]
  reg  flight_42; // @[FIFOFixer.scala 71:27]
  reg  flight_43; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_10; // @[Reg.scala 16:16]
  wire  stalls_10 = stalls_a_sel_10 & a_first & (flight_40 | flight_41 | flight_42 | flight_43) & (a_noDomain |
    stalls_id_10 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_11 = auto_in_a_bits_source[5:2] == 4'hb; // @[Parameters.scala 54:32]
  reg  flight_44; // @[FIFOFixer.scala 71:27]
  reg  flight_45; // @[FIFOFixer.scala 71:27]
  reg  flight_46; // @[FIFOFixer.scala 71:27]
  reg  flight_47; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_11; // @[Reg.scala 16:16]
  wire  stalls_11 = stalls_a_sel_11 & a_first & (flight_44 | flight_45 | flight_46 | flight_47) & (a_noDomain |
    stalls_id_11 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_12 = auto_in_a_bits_source[5:2] == 4'hc; // @[Parameters.scala 54:32]
  reg  flight_48; // @[FIFOFixer.scala 71:27]
  reg  flight_49; // @[FIFOFixer.scala 71:27]
  reg  flight_50; // @[FIFOFixer.scala 71:27]
  reg  flight_51; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_12; // @[Reg.scala 16:16]
  wire  stalls_12 = stalls_a_sel_12 & a_first & (flight_48 | flight_49 | flight_50 | flight_51) & (a_noDomain |
    stalls_id_12 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_13 = auto_in_a_bits_source[5:2] == 4'hd; // @[Parameters.scala 54:32]
  reg  flight_52; // @[FIFOFixer.scala 71:27]
  reg  flight_53; // @[FIFOFixer.scala 71:27]
  reg  flight_54; // @[FIFOFixer.scala 71:27]
  reg  flight_55; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_13; // @[Reg.scala 16:16]
  wire  stalls_13 = stalls_a_sel_13 & a_first & (flight_52 | flight_53 | flight_54 | flight_55) & (a_noDomain |
    stalls_id_13 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_14 = auto_in_a_bits_source[5:2] == 4'he; // @[Parameters.scala 54:32]
  reg  flight_56; // @[FIFOFixer.scala 71:27]
  reg  flight_57; // @[FIFOFixer.scala 71:27]
  reg  flight_58; // @[FIFOFixer.scala 71:27]
  reg  flight_59; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_14; // @[Reg.scala 16:16]
  wire  stalls_14 = stalls_a_sel_14 & a_first & (flight_56 | flight_57 | flight_58 | flight_59) & (a_noDomain |
    stalls_id_14 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stalls_a_sel_15 = auto_in_a_bits_source[5:2] == 4'hf; // @[Parameters.scala 54:32]
  reg  flight_60; // @[FIFOFixer.scala 71:27]
  reg  flight_61; // @[FIFOFixer.scala 71:27]
  reg  flight_62; // @[FIFOFixer.scala 71:27]
  reg  flight_63; // @[FIFOFixer.scala 71:27]
  reg  stalls_id_15; // @[Reg.scala 16:16]
  wire  stalls_15 = stalls_a_sel_15 & a_first & (flight_60 | flight_61 | flight_62 | flight_63) & (a_noDomain |
    stalls_id_15 != a_id); // @[FIFOFixer.scala 80:50]
  wire  stall = stalls_0 | stalls_1 | stalls_2 | stalls_3 | stalls_4 | stalls_5 | stalls_6 | stalls_7 | stalls_8 |
    stalls_9 | stalls_10 | stalls_11 | stalls_12 | stalls_13 | stalls_14 | stalls_15; // @[FIFOFixer.scala 83:49]
  wire  _bundleIn_0_a_ready_T = ~stall; // @[FIFOFixer.scala 88:50]
  wire  bundleIn_0_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  wire  _a_first_T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _a_first_beats1_decode_T_1 = 27'hfff << auto_in_a_bits_size; // @[package.scala 234:77]
  wire [11:0] _a_first_beats1_decode_T_3 = ~_a_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] a_first_beats1_decode = _a_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28]
  wire  _d_first_T = auto_in_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28]
  wire  d_first_first = d_first_counter == 9'h0; // @[Edges.scala 230:25]
  wire  d_first = d_first_first & auto_out_d_bits_opcode != 3'h6; // @[FIFOFixer.scala 67:42]
  wire  _GEN_66 = a_first & _a_first_T ? 6'h0 == auto_in_a_bits_source | flight_0 : flight_0; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_67 = a_first & _a_first_T ? 6'h1 == auto_in_a_bits_source | flight_1 : flight_1; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_68 = a_first & _a_first_T ? 6'h2 == auto_in_a_bits_source | flight_2 : flight_2; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_69 = a_first & _a_first_T ? 6'h3 == auto_in_a_bits_source | flight_3 : flight_3; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_70 = a_first & _a_first_T ? 6'h4 == auto_in_a_bits_source | flight_4 : flight_4; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_71 = a_first & _a_first_T ? 6'h5 == auto_in_a_bits_source | flight_5 : flight_5; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_72 = a_first & _a_first_T ? 6'h6 == auto_in_a_bits_source | flight_6 : flight_6; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_73 = a_first & _a_first_T ? 6'h7 == auto_in_a_bits_source | flight_7 : flight_7; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_74 = a_first & _a_first_T ? 6'h8 == auto_in_a_bits_source | flight_8 : flight_8; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_75 = a_first & _a_first_T ? 6'h9 == auto_in_a_bits_source | flight_9 : flight_9; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_76 = a_first & _a_first_T ? 6'ha == auto_in_a_bits_source | flight_10 : flight_10; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_77 = a_first & _a_first_T ? 6'hb == auto_in_a_bits_source | flight_11 : flight_11; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_78 = a_first & _a_first_T ? 6'hc == auto_in_a_bits_source | flight_12 : flight_12; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_79 = a_first & _a_first_T ? 6'hd == auto_in_a_bits_source | flight_13 : flight_13; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_80 = a_first & _a_first_T ? 6'he == auto_in_a_bits_source | flight_14 : flight_14; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_81 = a_first & _a_first_T ? 6'hf == auto_in_a_bits_source | flight_15 : flight_15; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_82 = a_first & _a_first_T ? 6'h10 == auto_in_a_bits_source | flight_16 : flight_16; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_83 = a_first & _a_first_T ? 6'h11 == auto_in_a_bits_source | flight_17 : flight_17; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_84 = a_first & _a_first_T ? 6'h12 == auto_in_a_bits_source | flight_18 : flight_18; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_85 = a_first & _a_first_T ? 6'h13 == auto_in_a_bits_source | flight_19 : flight_19; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_86 = a_first & _a_first_T ? 6'h14 == auto_in_a_bits_source | flight_20 : flight_20; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_87 = a_first & _a_first_T ? 6'h15 == auto_in_a_bits_source | flight_21 : flight_21; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_88 = a_first & _a_first_T ? 6'h16 == auto_in_a_bits_source | flight_22 : flight_22; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_89 = a_first & _a_first_T ? 6'h17 == auto_in_a_bits_source | flight_23 : flight_23; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_90 = a_first & _a_first_T ? 6'h18 == auto_in_a_bits_source | flight_24 : flight_24; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_91 = a_first & _a_first_T ? 6'h19 == auto_in_a_bits_source | flight_25 : flight_25; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_92 = a_first & _a_first_T ? 6'h1a == auto_in_a_bits_source | flight_26 : flight_26; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_93 = a_first & _a_first_T ? 6'h1b == auto_in_a_bits_source | flight_27 : flight_27; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_94 = a_first & _a_first_T ? 6'h1c == auto_in_a_bits_source | flight_28 : flight_28; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_95 = a_first & _a_first_T ? 6'h1d == auto_in_a_bits_source | flight_29 : flight_29; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_96 = a_first & _a_first_T ? 6'h1e == auto_in_a_bits_source | flight_30 : flight_30; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_97 = a_first & _a_first_T ? 6'h1f == auto_in_a_bits_source | flight_31 : flight_31; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_98 = a_first & _a_first_T ? 6'h20 == auto_in_a_bits_source | flight_32 : flight_32; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_99 = a_first & _a_first_T ? 6'h21 == auto_in_a_bits_source | flight_33 : flight_33; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_100 = a_first & _a_first_T ? 6'h22 == auto_in_a_bits_source | flight_34 : flight_34; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_101 = a_first & _a_first_T ? 6'h23 == auto_in_a_bits_source | flight_35 : flight_35; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_102 = a_first & _a_first_T ? 6'h24 == auto_in_a_bits_source | flight_36 : flight_36; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_103 = a_first & _a_first_T ? 6'h25 == auto_in_a_bits_source | flight_37 : flight_37; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_104 = a_first & _a_first_T ? 6'h26 == auto_in_a_bits_source | flight_38 : flight_38; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_105 = a_first & _a_first_T ? 6'h27 == auto_in_a_bits_source | flight_39 : flight_39; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_106 = a_first & _a_first_T ? 6'h28 == auto_in_a_bits_source | flight_40 : flight_40; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_107 = a_first & _a_first_T ? 6'h29 == auto_in_a_bits_source | flight_41 : flight_41; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_108 = a_first & _a_first_T ? 6'h2a == auto_in_a_bits_source | flight_42 : flight_42; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_109 = a_first & _a_first_T ? 6'h2b == auto_in_a_bits_source | flight_43 : flight_43; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_110 = a_first & _a_first_T ? 6'h2c == auto_in_a_bits_source | flight_44 : flight_44; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_111 = a_first & _a_first_T ? 6'h2d == auto_in_a_bits_source | flight_45 : flight_45; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_112 = a_first & _a_first_T ? 6'h2e == auto_in_a_bits_source | flight_46 : flight_46; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_113 = a_first & _a_first_T ? 6'h2f == auto_in_a_bits_source | flight_47 : flight_47; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_114 = a_first & _a_first_T ? 6'h30 == auto_in_a_bits_source | flight_48 : flight_48; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_115 = a_first & _a_first_T ? 6'h31 == auto_in_a_bits_source | flight_49 : flight_49; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_116 = a_first & _a_first_T ? 6'h32 == auto_in_a_bits_source | flight_50 : flight_50; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_117 = a_first & _a_first_T ? 6'h33 == auto_in_a_bits_source | flight_51 : flight_51; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_118 = a_first & _a_first_T ? 6'h34 == auto_in_a_bits_source | flight_52 : flight_52; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_119 = a_first & _a_first_T ? 6'h35 == auto_in_a_bits_source | flight_53 : flight_53; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_120 = a_first & _a_first_T ? 6'h36 == auto_in_a_bits_source | flight_54 : flight_54; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_121 = a_first & _a_first_T ? 6'h37 == auto_in_a_bits_source | flight_55 : flight_55; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_122 = a_first & _a_first_T ? 6'h38 == auto_in_a_bits_source | flight_56 : flight_56; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_123 = a_first & _a_first_T ? 6'h39 == auto_in_a_bits_source | flight_57 : flight_57; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_124 = a_first & _a_first_T ? 6'h3a == auto_in_a_bits_source | flight_58 : flight_58; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_125 = a_first & _a_first_T ? 6'h3b == auto_in_a_bits_source | flight_59 : flight_59; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_126 = a_first & _a_first_T ? 6'h3c == auto_in_a_bits_source | flight_60 : flight_60; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_127 = a_first & _a_first_T ? 6'h3d == auto_in_a_bits_source | flight_61 : flight_61; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_128 = a_first & _a_first_T ? 6'h3e == auto_in_a_bits_source | flight_62 : flight_62; // @[FIFOFixer.scala 71:27 72:37]
  wire  _GEN_129 = a_first & _a_first_T ? 6'h3f == auto_in_a_bits_source | flight_63 : flight_63; // @[FIFOFixer.scala 71:27 72:37]
  wire  _stalls_id_T_1 = _a_first_T & stalls_a_sel; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_5 = _a_first_T & stalls_a_sel_1; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_9 = _a_first_T & stalls_a_sel_2; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_13 = _a_first_T & stalls_a_sel_3; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_17 = _a_first_T & stalls_a_sel_4; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_21 = _a_first_T & stalls_a_sel_5; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_25 = _a_first_T & stalls_a_sel_6; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_29 = _a_first_T & stalls_a_sel_7; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_33 = _a_first_T & stalls_a_sel_8; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_37 = _a_first_T & stalls_a_sel_9; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_41 = _a_first_T & stalls_a_sel_10; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_45 = _a_first_T & stalls_a_sel_11; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_49 = _a_first_T & stalls_a_sel_12; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_53 = _a_first_T & stalls_a_sel_13; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_57 = _a_first_T & stalls_a_sel_14; // @[FIFOFixer.scala 77:49]
  wire  _stalls_id_T_61 = _a_first_T & stalls_a_sel_15; // @[FIFOFixer.scala 77:49]
  reg [16:0] TLFIFOFixer_5_covState; // @[Register tracking TLFIFOFixer_5 state]
  reg  TLFIFOFixer_5_covMap [0:131071]; // @[Coverage map for TLFIFOFixer_5]
  wire  TLFIFOFixer_5_covMap_read_en; // @[Coverage map for TLFIFOFixer_5]
  wire [16:0] TLFIFOFixer_5_covMap_read_addr; // @[Coverage map for TLFIFOFixer_5]
  wire  TLFIFOFixer_5_covMap_read_data; // @[Coverage map for TLFIFOFixer_5]
  wire  TLFIFOFixer_5_covMap_write_data; // @[Coverage map for TLFIFOFixer_5]
  wire [16:0] TLFIFOFixer_5_covMap_write_addr; // @[Coverage map for TLFIFOFixer_5]
  wire  TLFIFOFixer_5_covMap_write_mask; // @[Coverage map for TLFIFOFixer_5]
  wire  TLFIFOFixer_5_covMap_write_en; // @[Coverage map for TLFIFOFixer_5]
  reg [29:0] TLFIFOFixer_5_covSum; // @[Sum of coverage map]
  wire  stalls_id_8_shl;
  wire [16:0] stalls_id_8_pad;
  wire [1:0] stalls_id_7_shl;
  wire [16:0] stalls_id_7_pad;
  wire [2:0] stalls_id_shl;
  wire [16:0] stalls_id_pad;
  wire [3:0] stalls_id_6_shl;
  wire [16:0] stalls_id_6_pad;
  wire [4:0] stalls_id_15_shl;
  wire [16:0] stalls_id_15_pad;
  wire [5:0] stalls_id_9_shl;
  wire [16:0] stalls_id_9_pad;
  wire [6:0] stalls_id_5_shl;
  wire [16:0] stalls_id_5_pad;
  wire [7:0] stalls_id_2_shl;
  wire [16:0] stalls_id_2_pad;
  wire [8:0] stalls_id_3_shl;
  wire [16:0] stalls_id_3_pad;
  wire [9:0] stalls_id_12_shl;
  wire [16:0] stalls_id_12_pad;
  wire [10:0] stalls_id_11_shl;
  wire [16:0] stalls_id_11_pad;
  wire [11:0] stalls_id_13_shl;
  wire [16:0] stalls_id_13_pad;
  wire [12:0] stalls_id_4_shl;
  wire [16:0] stalls_id_4_pad;
  wire [13:0] stalls_id_1_shl;
  wire [16:0] stalls_id_1_pad;
  wire [14:0] stalls_id_10_shl;
  wire [16:0] stalls_id_10_pad;
  wire [15:0] stalls_id_14_shl;
  wire [16:0] stalls_id_14_pad;
  wire [16:0] flight_41_shl;
  wire [16:0] flight_41_pad;
  wire [16:0] flight_53_shl;
  wire [16:0] flight_53_pad;
  wire [16:0] flight_1_shl;
  wire [16:0] flight_1_pad;
  wire [16:0] flight_40_shl;
  wire [16:0] flight_40_pad;
  wire [16:0] flight_23_shl;
  wire [16:0] flight_23_pad;
  wire [16:0] flight_34_shl;
  wire [16:0] flight_34_pad;
  wire [16:0] flight_47_shl;
  wire [16:0] flight_47_pad;
  wire [16:0] flight_56_shl;
  wire [16:0] flight_56_pad;
  wire [16:0] flight_20_shl;
  wire [16:0] flight_20_pad;
  wire [16:0] flight_60_shl;
  wire [16:0] flight_60_pad;
  wire [16:0] flight_49_shl;
  wire [16:0] flight_49_pad;
  wire [16:0] flight_12_shl;
  wire [16:0] flight_12_pad;
  wire [16:0] flight_8_shl;
  wire [16:0] flight_8_pad;
  wire [16:0] flight_9_shl;
  wire [16:0] flight_9_pad;
  wire [16:0] flight_57_shl;
  wire [16:0] flight_57_pad;
  wire [16:0] flight_48_shl;
  wire [16:0] flight_48_pad;
  wire [16:0] flight_10_shl;
  wire [16:0] flight_10_pad;
  wire [16:0] flight_32_shl;
  wire [16:0] flight_32_pad;
  wire [16:0] flight_61_shl;
  wire [16:0] flight_61_pad;
  wire [16:0] flight_5_shl;
  wire [16:0] flight_5_pad;
  wire [16:0] flight_39_shl;
  wire [16:0] flight_39_pad;
  wire [16:0] flight_19_shl;
  wire [16:0] flight_19_pad;
  wire [16:0] flight_58_shl;
  wire [16:0] flight_58_pad;
  wire [16:0] flight_21_shl;
  wire [16:0] flight_21_pad;
  wire [16:0] flight_62_shl;
  wire [16:0] flight_62_pad;
  wire [16:0] flight_15_shl;
  wire [16:0] flight_15_pad;
  wire [16:0] flight_14_shl;
  wire [16:0] flight_14_pad;
  wire [16:0] flight_51_shl;
  wire [16:0] flight_51_pad;
  wire [16:0] flight_37_shl;
  wire [16:0] flight_37_pad;
  wire [16:0] flight_13_shl;
  wire [16:0] flight_13_pad;
  wire [16:0] flight_46_shl;
  wire [16:0] flight_46_pad;
  wire [16:0] flight_16_shl;
  wire [16:0] flight_16_pad;
  wire [16:0] flight_7_shl;
  wire [16:0] flight_7_pad;
  wire [16:0] flight_0_shl;
  wire [16:0] flight_0_pad;
  wire [16:0] flight_38_shl;
  wire [16:0] flight_38_pad;
  wire [16:0] flight_30_shl;
  wire [16:0] flight_30_pad;
  wire [16:0] flight_22_shl;
  wire [16:0] flight_22_pad;
  wire [16:0] flight_59_shl;
  wire [16:0] flight_59_pad;
  wire [16:0] flight_55_shl;
  wire [16:0] flight_55_pad;
  wire [16:0] flight_45_shl;
  wire [16:0] flight_45_pad;
  wire [16:0] flight_11_shl;
  wire [16:0] flight_11_pad;
  wire [16:0] flight_6_shl;
  wire [16:0] flight_6_pad;
  wire [16:0] flight_31_shl;
  wire [16:0] flight_31_pad;
  wire [16:0] flight_3_shl;
  wire [16:0] flight_3_pad;
  wire [16:0] flight_42_shl;
  wire [16:0] flight_42_pad;
  wire [16:0] flight_25_shl;
  wire [16:0] flight_25_pad;
  wire [16:0] flight_17_shl;
  wire [16:0] flight_17_pad;
  wire [16:0] flight_36_shl;
  wire [16:0] flight_36_pad;
  wire [16:0] flight_2_shl;
  wire [16:0] flight_2_pad;
  wire [16:0] flight_29_shl;
  wire [16:0] flight_29_pad;
  wire [16:0] flight_27_shl;
  wire [16:0] flight_27_pad;
  wire [16:0] flight_33_shl;
  wire [16:0] flight_33_pad;
  wire [16:0] flight_35_shl;
  wire [16:0] flight_35_pad;
  wire [16:0] flight_4_shl;
  wire [16:0] flight_4_pad;
  wire [16:0] flight_28_shl;
  wire [16:0] flight_28_pad;
  wire [16:0] flight_18_shl;
  wire [16:0] flight_18_pad;
  wire [16:0] flight_63_shl;
  wire [16:0] flight_63_pad;
  wire [16:0] flight_54_shl;
  wire [16:0] flight_54_pad;
  wire [16:0] flight_50_shl;
  wire [16:0] flight_50_pad;
  wire [16:0] flight_44_shl;
  wire [16:0] flight_44_pad;
  wire [16:0] flight_43_shl;
  wire [16:0] flight_43_pad;
  wire [16:0] flight_52_shl;
  wire [16:0] flight_52_pad;
  wire [16:0] flight_26_shl;
  wire [16:0] flight_26_pad;
  wire [16:0] flight_24_shl;
  wire [16:0] flight_24_pad;
  wire [16:0] TLFIFOFixer_5_xor31;
  wire [16:0] TLFIFOFixer_5_xor66;
  wire [16:0] TLFIFOFixer_5_xor32;
  wire [16:0] TLFIFOFixer_5_xor15;
  wire [16:0] TLFIFOFixer_5_xor33;
  wire [16:0] TLFIFOFixer_5_xor70;
  wire [16:0] TLFIFOFixer_5_xor34;
  wire [16:0] TLFIFOFixer_5_xor16;
  wire [16:0] TLFIFOFixer_5_xor7;
  wire [16:0] TLFIFOFixer_5_xor35;
  wire [16:0] TLFIFOFixer_5_xor74;
  wire [16:0] TLFIFOFixer_5_xor36;
  wire [16:0] TLFIFOFixer_5_xor17;
  wire [16:0] TLFIFOFixer_5_xor37;
  wire [16:0] TLFIFOFixer_5_xor78;
  wire [16:0] TLFIFOFixer_5_xor38;
  wire [16:0] TLFIFOFixer_5_xor18;
  wire [16:0] TLFIFOFixer_5_xor8;
  wire [16:0] TLFIFOFixer_5_xor3;
  wire [16:0] TLFIFOFixer_5_xor39;
  wire [16:0] TLFIFOFixer_5_xor82;
  wire [16:0] TLFIFOFixer_5_xor40;
  wire [16:0] TLFIFOFixer_5_xor19;
  wire [16:0] TLFIFOFixer_5_xor41;
  wire [16:0] TLFIFOFixer_5_xor86;
  wire [16:0] TLFIFOFixer_5_xor42;
  wire [16:0] TLFIFOFixer_5_xor20;
  wire [16:0] TLFIFOFixer_5_xor9;
  wire [16:0] TLFIFOFixer_5_xor43;
  wire [16:0] TLFIFOFixer_5_xor90;
  wire [16:0] TLFIFOFixer_5_xor44;
  wire [16:0] TLFIFOFixer_5_xor21;
  wire [16:0] TLFIFOFixer_5_xor45;
  wire [16:0] TLFIFOFixer_5_xor94;
  wire [16:0] TLFIFOFixer_5_xor46;
  wire [16:0] TLFIFOFixer_5_xor22;
  wire [16:0] TLFIFOFixer_5_xor10;
  wire [16:0] TLFIFOFixer_5_xor4;
  wire [16:0] TLFIFOFixer_5_xor1;
  wire [16:0] TLFIFOFixer_5_xor47;
  wire [16:0] TLFIFOFixer_5_xor98;
  wire [16:0] TLFIFOFixer_5_xor48;
  wire [16:0] TLFIFOFixer_5_xor23;
  wire [16:0] TLFIFOFixer_5_xor49;
  wire [16:0] TLFIFOFixer_5_xor102;
  wire [16:0] TLFIFOFixer_5_xor50;
  wire [16:0] TLFIFOFixer_5_xor24;
  wire [16:0] TLFIFOFixer_5_xor11;
  wire [16:0] TLFIFOFixer_5_xor51;
  wire [16:0] TLFIFOFixer_5_xor106;
  wire [16:0] TLFIFOFixer_5_xor52;
  wire [16:0] TLFIFOFixer_5_xor25;
  wire [16:0] TLFIFOFixer_5_xor53;
  wire [16:0] TLFIFOFixer_5_xor110;
  wire [16:0] TLFIFOFixer_5_xor54;
  wire [16:0] TLFIFOFixer_5_xor26;
  wire [16:0] TLFIFOFixer_5_xor12;
  wire [16:0] TLFIFOFixer_5_xor5;
  wire [16:0] TLFIFOFixer_5_xor55;
  wire [16:0] TLFIFOFixer_5_xor114;
  wire [16:0] TLFIFOFixer_5_xor56;
  wire [16:0] TLFIFOFixer_5_xor27;
  wire [16:0] TLFIFOFixer_5_xor57;
  wire [16:0] TLFIFOFixer_5_xor118;
  wire [16:0] TLFIFOFixer_5_xor58;
  wire [16:0] TLFIFOFixer_5_xor28;
  wire [16:0] TLFIFOFixer_5_xor13;
  wire [16:0] TLFIFOFixer_5_xor59;
  wire [16:0] TLFIFOFixer_5_xor122;
  wire [16:0] TLFIFOFixer_5_xor60;
  wire [16:0] TLFIFOFixer_5_xor29;
  wire [16:0] TLFIFOFixer_5_xor61;
  wire [16:0] TLFIFOFixer_5_xor126;
  wire [16:0] TLFIFOFixer_5_xor62;
  wire [16:0] TLFIFOFixer_5_xor30;
  wire [16:0] TLFIFOFixer_5_xor14;
  wire [16:0] TLFIFOFixer_5_xor6;
  wire [16:0] TLFIFOFixer_5_xor2;
  wire [16:0] TLFIFOFixer_5_xor0;
  assign auto_in_a_ready = auto_out_a_ready & ~stall; // @[FIFOFixer.scala 88:33]
  assign auto_in_d_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_a_valid = auto_in_a_valid & _bundleIn_0_a_ready_T; // @[FIFOFixer.scala 87:33]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_bufferable = auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_modifiable = auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_readalloc = auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_writealloc = auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_privileged = auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_secure = auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_user_amba_prot_fetch = auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign TLFIFOFixer_5_covMap_read_en = 1'h1;
  assign TLFIFOFixer_5_covMap_read_addr = TLFIFOFixer_5_covState;
  assign TLFIFOFixer_5_covMap_read_data = TLFIFOFixer_5_covMap[TLFIFOFixer_5_covMap_read_addr]; // @[Coverage map for TLFIFOFixer_5]
  assign TLFIFOFixer_5_covMap_write_data = 1'h1;
  assign TLFIFOFixer_5_covMap_write_addr = TLFIFOFixer_5_covState;
  assign TLFIFOFixer_5_covMap_write_mask = 1'h1;
  assign TLFIFOFixer_5_covMap_write_en = ~metaReset;
  assign stalls_id_8_shl = stalls_id_8;
  assign stalls_id_8_pad = {16'h0,stalls_id_8_shl};
  assign stalls_id_7_shl = {stalls_id_7, 1'h0};
  assign stalls_id_7_pad = {15'h0,stalls_id_7_shl};
  assign stalls_id_shl = {stalls_id, 2'h0};
  assign stalls_id_pad = {14'h0,stalls_id_shl};
  assign stalls_id_6_shl = {stalls_id_6, 3'h0};
  assign stalls_id_6_pad = {13'h0,stalls_id_6_shl};
  assign stalls_id_15_shl = {stalls_id_15, 4'h0};
  assign stalls_id_15_pad = {12'h0,stalls_id_15_shl};
  assign stalls_id_9_shl = {stalls_id_9, 5'h0};
  assign stalls_id_9_pad = {11'h0,stalls_id_9_shl};
  assign stalls_id_5_shl = {stalls_id_5, 6'h0};
  assign stalls_id_5_pad = {10'h0,stalls_id_5_shl};
  assign stalls_id_2_shl = {stalls_id_2, 7'h0};
  assign stalls_id_2_pad = {9'h0,stalls_id_2_shl};
  assign stalls_id_3_shl = {stalls_id_3, 8'h0};
  assign stalls_id_3_pad = {8'h0,stalls_id_3_shl};
  assign stalls_id_12_shl = {stalls_id_12, 9'h0};
  assign stalls_id_12_pad = {7'h0,stalls_id_12_shl};
  assign stalls_id_11_shl = {stalls_id_11, 10'h0};
  assign stalls_id_11_pad = {6'h0,stalls_id_11_shl};
  assign stalls_id_13_shl = {stalls_id_13, 11'h0};
  assign stalls_id_13_pad = {5'h0,stalls_id_13_shl};
  assign stalls_id_4_shl = {stalls_id_4, 12'h0};
  assign stalls_id_4_pad = {4'h0,stalls_id_4_shl};
  assign stalls_id_1_shl = {stalls_id_1, 13'h0};
  assign stalls_id_1_pad = {3'h0,stalls_id_1_shl};
  assign stalls_id_10_shl = {stalls_id_10, 14'h0};
  assign stalls_id_10_pad = {2'h0,stalls_id_10_shl};
  assign stalls_id_14_shl = {stalls_id_14, 15'h0};
  assign stalls_id_14_pad = {1'h0,stalls_id_14_shl};
  assign flight_41_shl = {flight_41, 16'h0};
  assign flight_41_pad = flight_41_shl;
  assign flight_53_shl = {flight_53, 16'h0};
  assign flight_53_pad = flight_53_shl;
  assign flight_1_shl = {flight_1, 16'h0};
  assign flight_1_pad = flight_1_shl;
  assign flight_40_shl = {flight_40, 16'h0};
  assign flight_40_pad = flight_40_shl;
  assign flight_23_shl = {flight_23, 16'h0};
  assign flight_23_pad = flight_23_shl;
  assign flight_34_shl = {flight_34, 16'h0};
  assign flight_34_pad = flight_34_shl;
  assign flight_47_shl = {flight_47, 16'h0};
  assign flight_47_pad = flight_47_shl;
  assign flight_56_shl = {flight_56, 16'h0};
  assign flight_56_pad = flight_56_shl;
  assign flight_20_shl = {flight_20, 16'h0};
  assign flight_20_pad = flight_20_shl;
  assign flight_60_shl = {flight_60, 16'h0};
  assign flight_60_pad = flight_60_shl;
  assign flight_49_shl = {flight_49, 16'h0};
  assign flight_49_pad = flight_49_shl;
  assign flight_12_shl = {flight_12, 16'h0};
  assign flight_12_pad = flight_12_shl;
  assign flight_8_shl = {flight_8, 16'h0};
  assign flight_8_pad = flight_8_shl;
  assign flight_9_shl = {flight_9, 16'h0};
  assign flight_9_pad = flight_9_shl;
  assign flight_57_shl = {flight_57, 16'h0};
  assign flight_57_pad = flight_57_shl;
  assign flight_48_shl = {flight_48, 16'h0};
  assign flight_48_pad = flight_48_shl;
  assign flight_10_shl = {flight_10, 16'h0};
  assign flight_10_pad = flight_10_shl;
  assign flight_32_shl = {flight_32, 16'h0};
  assign flight_32_pad = flight_32_shl;
  assign flight_61_shl = {flight_61, 16'h0};
  assign flight_61_pad = flight_61_shl;
  assign flight_5_shl = {flight_5, 16'h0};
  assign flight_5_pad = flight_5_shl;
  assign flight_39_shl = {flight_39, 16'h0};
  assign flight_39_pad = flight_39_shl;
  assign flight_19_shl = {flight_19, 16'h0};
  assign flight_19_pad = flight_19_shl;
  assign flight_58_shl = {flight_58, 16'h0};
  assign flight_58_pad = flight_58_shl;
  assign flight_21_shl = {flight_21, 16'h0};
  assign flight_21_pad = flight_21_shl;
  assign flight_62_shl = {flight_62, 16'h0};
  assign flight_62_pad = flight_62_shl;
  assign flight_15_shl = {flight_15, 16'h0};
  assign flight_15_pad = flight_15_shl;
  assign flight_14_shl = {flight_14, 16'h0};
  assign flight_14_pad = flight_14_shl;
  assign flight_51_shl = {flight_51, 16'h0};
  assign flight_51_pad = flight_51_shl;
  assign flight_37_shl = {flight_37, 16'h0};
  assign flight_37_pad = flight_37_shl;
  assign flight_13_shl = {flight_13, 16'h0};
  assign flight_13_pad = flight_13_shl;
  assign flight_46_shl = {flight_46, 16'h0};
  assign flight_46_pad = flight_46_shl;
  assign flight_16_shl = {flight_16, 16'h0};
  assign flight_16_pad = flight_16_shl;
  assign flight_7_shl = {flight_7, 16'h0};
  assign flight_7_pad = flight_7_shl;
  assign flight_0_shl = {flight_0, 16'h0};
  assign flight_0_pad = flight_0_shl;
  assign flight_38_shl = {flight_38, 16'h0};
  assign flight_38_pad = flight_38_shl;
  assign flight_30_shl = {flight_30, 16'h0};
  assign flight_30_pad = flight_30_shl;
  assign flight_22_shl = {flight_22, 16'h0};
  assign flight_22_pad = flight_22_shl;
  assign flight_59_shl = {flight_59, 16'h0};
  assign flight_59_pad = flight_59_shl;
  assign flight_55_shl = {flight_55, 16'h0};
  assign flight_55_pad = flight_55_shl;
  assign flight_45_shl = {flight_45, 16'h0};
  assign flight_45_pad = flight_45_shl;
  assign flight_11_shl = {flight_11, 16'h0};
  assign flight_11_pad = flight_11_shl;
  assign flight_6_shl = {flight_6, 16'h0};
  assign flight_6_pad = flight_6_shl;
  assign flight_31_shl = {flight_31, 16'h0};
  assign flight_31_pad = flight_31_shl;
  assign flight_3_shl = {flight_3, 16'h0};
  assign flight_3_pad = flight_3_shl;
  assign flight_42_shl = {flight_42, 16'h0};
  assign flight_42_pad = flight_42_shl;
  assign flight_25_shl = {flight_25, 16'h0};
  assign flight_25_pad = flight_25_shl;
  assign flight_17_shl = {flight_17, 16'h0};
  assign flight_17_pad = flight_17_shl;
  assign flight_36_shl = {flight_36, 16'h0};
  assign flight_36_pad = flight_36_shl;
  assign flight_2_shl = {flight_2, 16'h0};
  assign flight_2_pad = flight_2_shl;
  assign flight_29_shl = {flight_29, 16'h0};
  assign flight_29_pad = flight_29_shl;
  assign flight_27_shl = {flight_27, 16'h0};
  assign flight_27_pad = flight_27_shl;
  assign flight_33_shl = {flight_33, 16'h0};
  assign flight_33_pad = flight_33_shl;
  assign flight_35_shl = {flight_35, 16'h0};
  assign flight_35_pad = flight_35_shl;
  assign flight_4_shl = {flight_4, 16'h0};
  assign flight_4_pad = flight_4_shl;
  assign flight_28_shl = {flight_28, 16'h0};
  assign flight_28_pad = flight_28_shl;
  assign flight_18_shl = {flight_18, 16'h0};
  assign flight_18_pad = flight_18_shl;
  assign flight_63_shl = {flight_63, 16'h0};
  assign flight_63_pad = flight_63_shl;
  assign flight_54_shl = {flight_54, 16'h0};
  assign flight_54_pad = flight_54_shl;
  assign flight_50_shl = {flight_50, 16'h0};
  assign flight_50_pad = flight_50_shl;
  assign flight_44_shl = {flight_44, 16'h0};
  assign flight_44_pad = flight_44_shl;
  assign flight_43_shl = {flight_43, 16'h0};
  assign flight_43_pad = flight_43_shl;
  assign flight_52_shl = {flight_52, 16'h0};
  assign flight_52_pad = flight_52_shl;
  assign flight_26_shl = {flight_26, 16'h0};
  assign flight_26_pad = flight_26_shl;
  assign flight_24_shl = {flight_24, 16'h0};
  assign flight_24_pad = flight_24_shl;
  assign TLFIFOFixer_5_xor31 = stalls_id_8_pad ^ stalls_id_7_pad;
  assign TLFIFOFixer_5_xor66 = stalls_id_6_pad ^ stalls_id_15_pad;
  assign TLFIFOFixer_5_xor32 = stalls_id_pad ^ TLFIFOFixer_5_xor66;
  assign TLFIFOFixer_5_xor15 = TLFIFOFixer_5_xor31 ^ TLFIFOFixer_5_xor32;
  assign TLFIFOFixer_5_xor33 = stalls_id_9_pad ^ stalls_id_5_pad;
  assign TLFIFOFixer_5_xor70 = stalls_id_3_pad ^ stalls_id_12_pad;
  assign TLFIFOFixer_5_xor34 = stalls_id_2_pad ^ TLFIFOFixer_5_xor70;
  assign TLFIFOFixer_5_xor16 = TLFIFOFixer_5_xor33 ^ TLFIFOFixer_5_xor34;
  assign TLFIFOFixer_5_xor7 = TLFIFOFixer_5_xor15 ^ TLFIFOFixer_5_xor16;
  assign TLFIFOFixer_5_xor35 = stalls_id_11_pad ^ stalls_id_13_pad;
  assign TLFIFOFixer_5_xor74 = stalls_id_1_pad ^ stalls_id_10_pad;
  assign TLFIFOFixer_5_xor36 = stalls_id_4_pad ^ TLFIFOFixer_5_xor74;
  assign TLFIFOFixer_5_xor17 = TLFIFOFixer_5_xor35 ^ TLFIFOFixer_5_xor36;
  assign TLFIFOFixer_5_xor37 = stalls_id_14_pad ^ flight_41_pad;
  assign TLFIFOFixer_5_xor78 = flight_1_pad ^ flight_40_pad;
  assign TLFIFOFixer_5_xor38 = flight_53_pad ^ TLFIFOFixer_5_xor78;
  assign TLFIFOFixer_5_xor18 = TLFIFOFixer_5_xor37 ^ TLFIFOFixer_5_xor38;
  assign TLFIFOFixer_5_xor8 = TLFIFOFixer_5_xor17 ^ TLFIFOFixer_5_xor18;
  assign TLFIFOFixer_5_xor3 = TLFIFOFixer_5_xor7 ^ TLFIFOFixer_5_xor8;
  assign TLFIFOFixer_5_xor39 = flight_23_pad ^ flight_34_pad;
  assign TLFIFOFixer_5_xor82 = flight_56_pad ^ flight_20_pad;
  assign TLFIFOFixer_5_xor40 = flight_47_pad ^ TLFIFOFixer_5_xor82;
  assign TLFIFOFixer_5_xor19 = TLFIFOFixer_5_xor39 ^ TLFIFOFixer_5_xor40;
  assign TLFIFOFixer_5_xor41 = flight_60_pad ^ flight_49_pad;
  assign TLFIFOFixer_5_xor86 = flight_8_pad ^ flight_9_pad;
  assign TLFIFOFixer_5_xor42 = flight_12_pad ^ TLFIFOFixer_5_xor86;
  assign TLFIFOFixer_5_xor20 = TLFIFOFixer_5_xor41 ^ TLFIFOFixer_5_xor42;
  assign TLFIFOFixer_5_xor9 = TLFIFOFixer_5_xor19 ^ TLFIFOFixer_5_xor20;
  assign TLFIFOFixer_5_xor43 = flight_57_pad ^ flight_48_pad;
  assign TLFIFOFixer_5_xor90 = flight_32_pad ^ flight_61_pad;
  assign TLFIFOFixer_5_xor44 = flight_10_pad ^ TLFIFOFixer_5_xor90;
  assign TLFIFOFixer_5_xor21 = TLFIFOFixer_5_xor43 ^ TLFIFOFixer_5_xor44;
  assign TLFIFOFixer_5_xor45 = flight_5_pad ^ flight_39_pad;
  assign TLFIFOFixer_5_xor94 = flight_58_pad ^ flight_21_pad;
  assign TLFIFOFixer_5_xor46 = flight_19_pad ^ TLFIFOFixer_5_xor94;
  assign TLFIFOFixer_5_xor22 = TLFIFOFixer_5_xor45 ^ TLFIFOFixer_5_xor46;
  assign TLFIFOFixer_5_xor10 = TLFIFOFixer_5_xor21 ^ TLFIFOFixer_5_xor22;
  assign TLFIFOFixer_5_xor4 = TLFIFOFixer_5_xor9 ^ TLFIFOFixer_5_xor10;
  assign TLFIFOFixer_5_xor1 = TLFIFOFixer_5_xor3 ^ TLFIFOFixer_5_xor4;
  assign TLFIFOFixer_5_xor47 = flight_62_pad ^ flight_15_pad;
  assign TLFIFOFixer_5_xor98 = flight_51_pad ^ flight_37_pad;
  assign TLFIFOFixer_5_xor48 = flight_14_pad ^ TLFIFOFixer_5_xor98;
  assign TLFIFOFixer_5_xor23 = TLFIFOFixer_5_xor47 ^ TLFIFOFixer_5_xor48;
  assign TLFIFOFixer_5_xor49 = flight_13_pad ^ flight_46_pad;
  assign TLFIFOFixer_5_xor102 = flight_7_pad ^ flight_0_pad;
  assign TLFIFOFixer_5_xor50 = flight_16_pad ^ TLFIFOFixer_5_xor102;
  assign TLFIFOFixer_5_xor24 = TLFIFOFixer_5_xor49 ^ TLFIFOFixer_5_xor50;
  assign TLFIFOFixer_5_xor11 = TLFIFOFixer_5_xor23 ^ TLFIFOFixer_5_xor24;
  assign TLFIFOFixer_5_xor51 = flight_38_pad ^ flight_30_pad;
  assign TLFIFOFixer_5_xor106 = flight_59_pad ^ flight_55_pad;
  assign TLFIFOFixer_5_xor52 = flight_22_pad ^ TLFIFOFixer_5_xor106;
  assign TLFIFOFixer_5_xor25 = TLFIFOFixer_5_xor51 ^ TLFIFOFixer_5_xor52;
  assign TLFIFOFixer_5_xor53 = flight_45_pad ^ flight_11_pad;
  assign TLFIFOFixer_5_xor110 = flight_31_pad ^ flight_3_pad;
  assign TLFIFOFixer_5_xor54 = flight_6_pad ^ TLFIFOFixer_5_xor110;
  assign TLFIFOFixer_5_xor26 = TLFIFOFixer_5_xor53 ^ TLFIFOFixer_5_xor54;
  assign TLFIFOFixer_5_xor12 = TLFIFOFixer_5_xor25 ^ TLFIFOFixer_5_xor26;
  assign TLFIFOFixer_5_xor5 = TLFIFOFixer_5_xor11 ^ TLFIFOFixer_5_xor12;
  assign TLFIFOFixer_5_xor55 = flight_42_pad ^ flight_25_pad;
  assign TLFIFOFixer_5_xor114 = flight_36_pad ^ flight_2_pad;
  assign TLFIFOFixer_5_xor56 = flight_17_pad ^ TLFIFOFixer_5_xor114;
  assign TLFIFOFixer_5_xor27 = TLFIFOFixer_5_xor55 ^ TLFIFOFixer_5_xor56;
  assign TLFIFOFixer_5_xor57 = flight_29_pad ^ flight_27_pad;
  assign TLFIFOFixer_5_xor118 = flight_35_pad ^ flight_4_pad;
  assign TLFIFOFixer_5_xor58 = flight_33_pad ^ TLFIFOFixer_5_xor118;
  assign TLFIFOFixer_5_xor28 = TLFIFOFixer_5_xor57 ^ TLFIFOFixer_5_xor58;
  assign TLFIFOFixer_5_xor13 = TLFIFOFixer_5_xor27 ^ TLFIFOFixer_5_xor28;
  assign TLFIFOFixer_5_xor59 = flight_28_pad ^ flight_18_pad;
  assign TLFIFOFixer_5_xor122 = flight_54_pad ^ flight_50_pad;
  assign TLFIFOFixer_5_xor60 = flight_63_pad ^ TLFIFOFixer_5_xor122;
  assign TLFIFOFixer_5_xor29 = TLFIFOFixer_5_xor59 ^ TLFIFOFixer_5_xor60;
  assign TLFIFOFixer_5_xor61 = flight_44_pad ^ flight_43_pad;
  assign TLFIFOFixer_5_xor126 = flight_26_pad ^ flight_24_pad;
  assign TLFIFOFixer_5_xor62 = flight_52_pad ^ TLFIFOFixer_5_xor126;
  assign TLFIFOFixer_5_xor30 = TLFIFOFixer_5_xor61 ^ TLFIFOFixer_5_xor62;
  assign TLFIFOFixer_5_xor14 = TLFIFOFixer_5_xor29 ^ TLFIFOFixer_5_xor30;
  assign TLFIFOFixer_5_xor6 = TLFIFOFixer_5_xor13 ^ TLFIFOFixer_5_xor14;
  assign TLFIFOFixer_5_xor2 = TLFIFOFixer_5_xor5 ^ TLFIFOFixer_5_xor6;
  assign TLFIFOFixer_5_xor0 = TLFIFOFixer_5_xor1 ^ TLFIFOFixer_5_xor2;
  assign io_covSum = TLFIFOFixer_5_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_a_first_T) begin
      if (a_first) begin
        if (a_first_beats1_opdata) begin
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_0 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h0 == auto_out_d_bits_source) begin
        flight_0 <= 1'h0;
      end else begin
        flight_0 <= _GEN_66;
      end
    end else begin
      flight_0 <= _GEN_66;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_1 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h1 == auto_out_d_bits_source) begin
        flight_1 <= 1'h0;
      end else begin
        flight_1 <= _GEN_67;
      end
    end else begin
      flight_1 <= _GEN_67;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_2 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h2 == auto_out_d_bits_source) begin
        flight_2 <= 1'h0;
      end else begin
        flight_2 <= _GEN_68;
      end
    end else begin
      flight_2 <= _GEN_68;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_3 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h3 == auto_out_d_bits_source) begin
        flight_3 <= 1'h0;
      end else begin
        flight_3 <= _GEN_69;
      end
    end else begin
      flight_3 <= _GEN_69;
    end
    if (_stalls_id_T_1) begin // @[Reg.scala 17:18]
      stalls_id <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_4 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h4 == auto_out_d_bits_source) begin
        flight_4 <= 1'h0;
      end else begin
        flight_4 <= _GEN_70;
      end
    end else begin
      flight_4 <= _GEN_70;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_5 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h5 == auto_out_d_bits_source) begin
        flight_5 <= 1'h0;
      end else begin
        flight_5 <= _GEN_71;
      end
    end else begin
      flight_5 <= _GEN_71;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_6 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h6 == auto_out_d_bits_source) begin
        flight_6 <= 1'h0;
      end else begin
        flight_6 <= _GEN_72;
      end
    end else begin
      flight_6 <= _GEN_72;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_7 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h7 == auto_out_d_bits_source) begin
        flight_7 <= 1'h0;
      end else begin
        flight_7 <= _GEN_73;
      end
    end else begin
      flight_7 <= _GEN_73;
    end
    if (_stalls_id_T_5) begin // @[Reg.scala 17:18]
      stalls_id_1 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_8 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h8 == auto_out_d_bits_source) begin
        flight_8 <= 1'h0;
      end else begin
        flight_8 <= _GEN_74;
      end
    end else begin
      flight_8 <= _GEN_74;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_9 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h9 == auto_out_d_bits_source) begin
        flight_9 <= 1'h0;
      end else begin
        flight_9 <= _GEN_75;
      end
    end else begin
      flight_9 <= _GEN_75;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_10 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'ha == auto_out_d_bits_source) begin
        flight_10 <= 1'h0;
      end else begin
        flight_10 <= _GEN_76;
      end
    end else begin
      flight_10 <= _GEN_76;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_11 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'hb == auto_out_d_bits_source) begin
        flight_11 <= 1'h0;
      end else begin
        flight_11 <= _GEN_77;
      end
    end else begin
      flight_11 <= _GEN_77;
    end
    if (_stalls_id_T_9) begin // @[Reg.scala 17:18]
      stalls_id_2 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_12 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'hc == auto_out_d_bits_source) begin
        flight_12 <= 1'h0;
      end else begin
        flight_12 <= _GEN_78;
      end
    end else begin
      flight_12 <= _GEN_78;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_13 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'hd == auto_out_d_bits_source) begin
        flight_13 <= 1'h0;
      end else begin
        flight_13 <= _GEN_79;
      end
    end else begin
      flight_13 <= _GEN_79;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_14 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'he == auto_out_d_bits_source) begin
        flight_14 <= 1'h0;
      end else begin
        flight_14 <= _GEN_80;
      end
    end else begin
      flight_14 <= _GEN_80;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_15 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'hf == auto_out_d_bits_source) begin
        flight_15 <= 1'h0;
      end else begin
        flight_15 <= _GEN_81;
      end
    end else begin
      flight_15 <= _GEN_81;
    end
    if (_stalls_id_T_13) begin // @[Reg.scala 17:18]
      stalls_id_3 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_16 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h10 == auto_out_d_bits_source) begin
        flight_16 <= 1'h0;
      end else begin
        flight_16 <= _GEN_82;
      end
    end else begin
      flight_16 <= _GEN_82;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_17 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h11 == auto_out_d_bits_source) begin
        flight_17 <= 1'h0;
      end else begin
        flight_17 <= _GEN_83;
      end
    end else begin
      flight_17 <= _GEN_83;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_18 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h12 == auto_out_d_bits_source) begin
        flight_18 <= 1'h0;
      end else begin
        flight_18 <= _GEN_84;
      end
    end else begin
      flight_18 <= _GEN_84;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_19 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h13 == auto_out_d_bits_source) begin
        flight_19 <= 1'h0;
      end else begin
        flight_19 <= _GEN_85;
      end
    end else begin
      flight_19 <= _GEN_85;
    end
    if (_stalls_id_T_17) begin // @[Reg.scala 17:18]
      stalls_id_4 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_20 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h14 == auto_out_d_bits_source) begin
        flight_20 <= 1'h0;
      end else begin
        flight_20 <= _GEN_86;
      end
    end else begin
      flight_20 <= _GEN_86;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_21 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h15 == auto_out_d_bits_source) begin
        flight_21 <= 1'h0;
      end else begin
        flight_21 <= _GEN_87;
      end
    end else begin
      flight_21 <= _GEN_87;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_22 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h16 == auto_out_d_bits_source) begin
        flight_22 <= 1'h0;
      end else begin
        flight_22 <= _GEN_88;
      end
    end else begin
      flight_22 <= _GEN_88;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_23 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h17 == auto_out_d_bits_source) begin
        flight_23 <= 1'h0;
      end else begin
        flight_23 <= _GEN_89;
      end
    end else begin
      flight_23 <= _GEN_89;
    end
    if (_stalls_id_T_21) begin // @[Reg.scala 17:18]
      stalls_id_5 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_24 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h18 == auto_out_d_bits_source) begin
        flight_24 <= 1'h0;
      end else begin
        flight_24 <= _GEN_90;
      end
    end else begin
      flight_24 <= _GEN_90;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_25 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h19 == auto_out_d_bits_source) begin
        flight_25 <= 1'h0;
      end else begin
        flight_25 <= _GEN_91;
      end
    end else begin
      flight_25 <= _GEN_91;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_26 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h1a == auto_out_d_bits_source) begin
        flight_26 <= 1'h0;
      end else begin
        flight_26 <= _GEN_92;
      end
    end else begin
      flight_26 <= _GEN_92;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_27 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h1b == auto_out_d_bits_source) begin
        flight_27 <= 1'h0;
      end else begin
        flight_27 <= _GEN_93;
      end
    end else begin
      flight_27 <= _GEN_93;
    end
    if (_stalls_id_T_25) begin // @[Reg.scala 17:18]
      stalls_id_6 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_28 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h1c == auto_out_d_bits_source) begin
        flight_28 <= 1'h0;
      end else begin
        flight_28 <= _GEN_94;
      end
    end else begin
      flight_28 <= _GEN_94;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_29 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h1d == auto_out_d_bits_source) begin
        flight_29 <= 1'h0;
      end else begin
        flight_29 <= _GEN_95;
      end
    end else begin
      flight_29 <= _GEN_95;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_30 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h1e == auto_out_d_bits_source) begin
        flight_30 <= 1'h0;
      end else begin
        flight_30 <= _GEN_96;
      end
    end else begin
      flight_30 <= _GEN_96;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_31 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h1f == auto_out_d_bits_source) begin
        flight_31 <= 1'h0;
      end else begin
        flight_31 <= _GEN_97;
      end
    end else begin
      flight_31 <= _GEN_97;
    end
    if (_stalls_id_T_29) begin // @[Reg.scala 17:18]
      stalls_id_7 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_32 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h20 == auto_out_d_bits_source) begin
        flight_32 <= 1'h0;
      end else begin
        flight_32 <= _GEN_98;
      end
    end else begin
      flight_32 <= _GEN_98;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_33 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h21 == auto_out_d_bits_source) begin
        flight_33 <= 1'h0;
      end else begin
        flight_33 <= _GEN_99;
      end
    end else begin
      flight_33 <= _GEN_99;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_34 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h22 == auto_out_d_bits_source) begin
        flight_34 <= 1'h0;
      end else begin
        flight_34 <= _GEN_100;
      end
    end else begin
      flight_34 <= _GEN_100;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_35 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h23 == auto_out_d_bits_source) begin
        flight_35 <= 1'h0;
      end else begin
        flight_35 <= _GEN_101;
      end
    end else begin
      flight_35 <= _GEN_101;
    end
    if (_stalls_id_T_33) begin // @[Reg.scala 17:18]
      stalls_id_8 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_36 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h24 == auto_out_d_bits_source) begin
        flight_36 <= 1'h0;
      end else begin
        flight_36 <= _GEN_102;
      end
    end else begin
      flight_36 <= _GEN_102;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_37 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h25 == auto_out_d_bits_source) begin
        flight_37 <= 1'h0;
      end else begin
        flight_37 <= _GEN_103;
      end
    end else begin
      flight_37 <= _GEN_103;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_38 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h26 == auto_out_d_bits_source) begin
        flight_38 <= 1'h0;
      end else begin
        flight_38 <= _GEN_104;
      end
    end else begin
      flight_38 <= _GEN_104;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_39 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h27 == auto_out_d_bits_source) begin
        flight_39 <= 1'h0;
      end else begin
        flight_39 <= _GEN_105;
      end
    end else begin
      flight_39 <= _GEN_105;
    end
    if (_stalls_id_T_37) begin // @[Reg.scala 17:18]
      stalls_id_9 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_40 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h28 == auto_out_d_bits_source) begin
        flight_40 <= 1'h0;
      end else begin
        flight_40 <= _GEN_106;
      end
    end else begin
      flight_40 <= _GEN_106;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_41 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h29 == auto_out_d_bits_source) begin
        flight_41 <= 1'h0;
      end else begin
        flight_41 <= _GEN_107;
      end
    end else begin
      flight_41 <= _GEN_107;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_42 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h2a == auto_out_d_bits_source) begin
        flight_42 <= 1'h0;
      end else begin
        flight_42 <= _GEN_108;
      end
    end else begin
      flight_42 <= _GEN_108;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_43 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h2b == auto_out_d_bits_source) begin
        flight_43 <= 1'h0;
      end else begin
        flight_43 <= _GEN_109;
      end
    end else begin
      flight_43 <= _GEN_109;
    end
    if (_stalls_id_T_41) begin // @[Reg.scala 17:18]
      stalls_id_10 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_44 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h2c == auto_out_d_bits_source) begin
        flight_44 <= 1'h0;
      end else begin
        flight_44 <= _GEN_110;
      end
    end else begin
      flight_44 <= _GEN_110;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_45 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h2d == auto_out_d_bits_source) begin
        flight_45 <= 1'h0;
      end else begin
        flight_45 <= _GEN_111;
      end
    end else begin
      flight_45 <= _GEN_111;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_46 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h2e == auto_out_d_bits_source) begin
        flight_46 <= 1'h0;
      end else begin
        flight_46 <= _GEN_112;
      end
    end else begin
      flight_46 <= _GEN_112;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_47 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h2f == auto_out_d_bits_source) begin
        flight_47 <= 1'h0;
      end else begin
        flight_47 <= _GEN_113;
      end
    end else begin
      flight_47 <= _GEN_113;
    end
    if (_stalls_id_T_45) begin // @[Reg.scala 17:18]
      stalls_id_11 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_48 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h30 == auto_out_d_bits_source) begin
        flight_48 <= 1'h0;
      end else begin
        flight_48 <= _GEN_114;
      end
    end else begin
      flight_48 <= _GEN_114;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_49 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h31 == auto_out_d_bits_source) begin
        flight_49 <= 1'h0;
      end else begin
        flight_49 <= _GEN_115;
      end
    end else begin
      flight_49 <= _GEN_115;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_50 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h32 == auto_out_d_bits_source) begin
        flight_50 <= 1'h0;
      end else begin
        flight_50 <= _GEN_116;
      end
    end else begin
      flight_50 <= _GEN_116;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_51 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h33 == auto_out_d_bits_source) begin
        flight_51 <= 1'h0;
      end else begin
        flight_51 <= _GEN_117;
      end
    end else begin
      flight_51 <= _GEN_117;
    end
    if (_stalls_id_T_49) begin // @[Reg.scala 17:18]
      stalls_id_12 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_52 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h34 == auto_out_d_bits_source) begin
        flight_52 <= 1'h0;
      end else begin
        flight_52 <= _GEN_118;
      end
    end else begin
      flight_52 <= _GEN_118;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_53 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h35 == auto_out_d_bits_source) begin
        flight_53 <= 1'h0;
      end else begin
        flight_53 <= _GEN_119;
      end
    end else begin
      flight_53 <= _GEN_119;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_54 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h36 == auto_out_d_bits_source) begin
        flight_54 <= 1'h0;
      end else begin
        flight_54 <= _GEN_120;
      end
    end else begin
      flight_54 <= _GEN_120;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_55 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h37 == auto_out_d_bits_source) begin
        flight_55 <= 1'h0;
      end else begin
        flight_55 <= _GEN_121;
      end
    end else begin
      flight_55 <= _GEN_121;
    end
    if (_stalls_id_T_53) begin // @[Reg.scala 17:18]
      stalls_id_13 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_56 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h38 == auto_out_d_bits_source) begin
        flight_56 <= 1'h0;
      end else begin
        flight_56 <= _GEN_122;
      end
    end else begin
      flight_56 <= _GEN_122;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_57 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h39 == auto_out_d_bits_source) begin
        flight_57 <= 1'h0;
      end else begin
        flight_57 <= _GEN_123;
      end
    end else begin
      flight_57 <= _GEN_123;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_58 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h3a == auto_out_d_bits_source) begin
        flight_58 <= 1'h0;
      end else begin
        flight_58 <= _GEN_124;
      end
    end else begin
      flight_58 <= _GEN_124;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_59 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h3b == auto_out_d_bits_source) begin
        flight_59 <= 1'h0;
      end else begin
        flight_59 <= _GEN_125;
      end
    end else begin
      flight_59 <= _GEN_125;
    end
    if (_stalls_id_T_57) begin // @[Reg.scala 17:18]
      stalls_id_14 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_60 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h3c == auto_out_d_bits_source) begin
        flight_60 <= 1'h0;
      end else begin
        flight_60 <= _GEN_126;
      end
    end else begin
      flight_60 <= _GEN_126;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_61 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h3d == auto_out_d_bits_source) begin
        flight_61 <= 1'h0;
      end else begin
        flight_61 <= _GEN_127;
      end
    end else begin
      flight_61 <= _GEN_127;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_62 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h3e == auto_out_d_bits_source) begin
        flight_62 <= 1'h0;
      end else begin
        flight_62 <= _GEN_128;
      end
    end else begin
      flight_62 <= _GEN_128;
    end
    if (reset) begin // @[FIFOFixer.scala 71:27]
      flight_63 <= 1'h0; // @[FIFOFixer.scala 71:27]
    end else if (d_first & _d_first_T) begin
      if (6'h3f == auto_out_d_bits_source) begin
        flight_63 <= 1'h0;
      end else begin
        flight_63 <= _GEN_129;
      end
    end else begin
      flight_63 <= _GEN_129;
    end
    if (_stalls_id_T_61) begin // @[Reg.scala 17:18]
      stalls_id_15 <= a_id; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_d_first_T) begin
      if (d_first_first) begin
        if (d_first_beats1_opdata) begin
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    TLFIFOFixer_5_covState <= TLFIFOFixer_5_xor0;
    if (TLFIFOFixer_5_covMap_write_en & TLFIFOFixer_5_covMap_write_mask) begin
      TLFIFOFixer_5_covMap[TLFIFOFixer_5_covMap_write_addr] <= TLFIFOFixer_5_covMap_write_data; // @[Coverage map for TLFIFOFixer_5]
    end
    if (!(TLFIFOFixer_5_covMap_read_data | metaReset)) begin
      TLFIFOFixer_5_covSum <= TLFIFOFixer_5_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_83 = {1{`RANDOM}};
  for (initvar = 0; initvar < 131072; initvar = initvar+1)
    TLFIFOFixer_5_covMap[initvar] = 0; //_83[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  flight_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  flight_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  flight_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  flight_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  stalls_id = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  flight_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  flight_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  flight_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  flight_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  stalls_id_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  flight_8 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  flight_9 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  flight_10 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  flight_11 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  stalls_id_2 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  flight_12 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  flight_13 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  flight_14 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  flight_15 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  stalls_id_3 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  flight_16 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  flight_17 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  flight_18 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  flight_19 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  stalls_id_4 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  flight_20 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  flight_21 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  flight_22 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  flight_23 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  stalls_id_5 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  flight_24 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  flight_25 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  flight_26 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  flight_27 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  stalls_id_6 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  flight_28 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  flight_29 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  flight_30 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  flight_31 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  stalls_id_7 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  flight_32 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  flight_33 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  flight_34 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  flight_35 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  stalls_id_8 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  flight_36 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  flight_37 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  flight_38 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  flight_39 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  stalls_id_9 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  flight_40 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  flight_41 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  flight_42 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  flight_43 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  stalls_id_10 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  flight_44 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  flight_45 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  flight_46 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  flight_47 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  stalls_id_11 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  flight_48 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  flight_49 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  flight_50 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  flight_51 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  stalls_id_12 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  flight_52 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  flight_53 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  flight_54 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  flight_55 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  stalls_id_13 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  flight_56 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  flight_57 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  flight_58 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  flight_59 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  stalls_id_14 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  flight_60 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  flight_61 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  flight_62 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  flight_63 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  stalls_id_15 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  d_first_counter = _RAND_81[8:0];
  _RAND_82 = {1{`RANDOM}};
  TLFIFOFixer_5_covState = 0; //_82[16:0];
  _RAND_84 = {1{`RANDOM}};
  TLFIFOFixer_5_covSum = 0; //_84[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_26(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_resp [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 259:95]
  reg  ram_last [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_12 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_12 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  reg  Queue_26_covState; // @[Register tracking Queue_26 state]
  reg  Queue_26_covMap [0:1]; // @[Coverage map for Queue_26]
  wire  Queue_26_covMap_read_en; // @[Coverage map for Queue_26]
  wire  Queue_26_covMap_read_addr; // @[Coverage map for Queue_26]
  wire  Queue_26_covMap_read_data; // @[Coverage map for Queue_26]
  wire  Queue_26_covMap_write_data; // @[Coverage map for Queue_26]
  wire  Queue_26_covMap_write_addr; // @[Coverage map for Queue_26]
  wire  Queue_26_covMap_write_mask; // @[Coverage map for Queue_26]
  wire  Queue_26_covMap_write_en; // @[Coverage map for Queue_26]
  reg [29:0] Queue_26_covSum; // @[Sum of coverage map]
  wire  maybe_full_shl;
  wire  maybe_full_pad;
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = 1'h0;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_12 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_resp = empty ? io_enq_bits_resp : ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_last = empty ? io_enq_bits_last : ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign Queue_26_covMap_read_en = 1'h1;
  assign Queue_26_covMap_read_addr = Queue_26_covState;
  assign Queue_26_covMap_read_data = Queue_26_covMap[Queue_26_covMap_read_addr]; // @[Coverage map for Queue_26]
  assign Queue_26_covMap_write_data = 1'h1;
  assign Queue_26_covMap_write_addr = Queue_26_covState;
  assign Queue_26_covMap_write_mask = 1'h1;
  assign Queue_26_covMap_write_en = ~metaReset;
  assign maybe_full_shl = maybe_full;
  assign maybe_full_pad = maybe_full_shl;
  assign io_covSum = Queue_26_covSum;
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
    Queue_26_covState <= maybe_full_pad;
    if (Queue_26_covMap_write_en & Queue_26_covMap_write_mask) begin
      Queue_26_covMap[Queue_26_covMap_write_addr] <= Queue_26_covMap_write_data; // @[Coverage map for Queue_26]
    end
    if (!(Queue_26_covMap_read_data | metaReset)) begin
      Queue_26_covSum <= Queue_26_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_3[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Queue_26_covMap[initvar] = 0; //_6[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  Queue_26_covState = 0; //_5[0:0];
  _RAND_7 = {1{`RANDOM}};
  Queue_26_covSum = 0; //_7[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_27(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [1:0]  io_enq_bits_resp,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [1:0]  io_deq_bits_resp,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_resp [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_resp_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_resp_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_10 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_10 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  reg  Queue_27_covState; // @[Register tracking Queue_27 state]
  reg  Queue_27_covMap [0:1]; // @[Coverage map for Queue_27]
  wire  Queue_27_covMap_read_en; // @[Coverage map for Queue_27]
  wire  Queue_27_covMap_read_addr; // @[Coverage map for Queue_27]
  wire  Queue_27_covMap_read_data; // @[Coverage map for Queue_27]
  wire  Queue_27_covMap_write_data; // @[Coverage map for Queue_27]
  wire  Queue_27_covMap_write_addr; // @[Coverage map for Queue_27]
  wire  Queue_27_covMap_write_mask; // @[Coverage map for Queue_27]
  wire  Queue_27_covMap_write_en; // @[Coverage map for Queue_27]
  reg [29:0] Queue_27_covSum; // @[Sum of coverage map]
  wire  maybe_full_shl;
  wire  maybe_full_pad;
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = 1'h0;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = empty ? _GEN_10 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_resp = empty ? io_enq_bits_resp : ram_resp_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign Queue_27_covMap_read_en = 1'h1;
  assign Queue_27_covMap_read_addr = Queue_27_covState;
  assign Queue_27_covMap_read_data = Queue_27_covMap[Queue_27_covMap_read_addr]; // @[Coverage map for Queue_27]
  assign Queue_27_covMap_write_data = 1'h1;
  assign Queue_27_covMap_write_addr = Queue_27_covState;
  assign Queue_27_covMap_write_mask = 1'h1;
  assign Queue_27_covMap_write_en = ~metaReset;
  assign maybe_full_shl = maybe_full;
  assign maybe_full_pad = maybe_full_shl;
  assign io_covSum = Queue_27_covSum;
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
    Queue_27_covState <= maybe_full_pad;
    if (Queue_27_covMap_write_en & Queue_27_covMap_write_mask) begin
      Queue_27_covMap[Queue_27_covMap_write_addr] <= Queue_27_covMap_write_data; // @[Coverage map for Queue_27]
    end
    if (!(Queue_27_covMap_read_data | metaReset)) begin
      Queue_27_covSum <= Queue_27_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = _RAND_1[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Queue_27_covMap[initvar] = 0; //_4[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  Queue_27_covState = 0; //_3[0:0];
  _RAND_5 = {1{`RANDOM}};
  Queue_27_covSum = 0; //_5[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4ToTL_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [3:0]  auto_out_a_bits_size,
  output [5:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output        auto_out_a_bits_user_amba_prot_bufferable,
  output        auto_out_a_bits_user_amba_prot_modifiable,
  output        auto_out_a_bits_user_amba_prot_readalloc,
  output        auto_out_a_bits_user_amba_prot_writealloc,
  output        auto_out_a_bits_user_amba_prot_privileged,
  output        auto_out_a_bits_user_amba_prot_secure,
  output        auto_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [3:0]  auto_out_d_bits_size,
  input  [5:0]  auto_out_d_bits_source,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_54;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_55;
`endif // RANDOMIZE_REG_INIT
  wire  deq_clock; // @[Decoupled.scala 361:21]
  wire  deq_reset; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] deq_io_enq_bits_id; // @[Decoupled.scala 361:21]
  wire [63:0] deq_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire [1:0] deq_io_enq_bits_resp; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_bits_last; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] deq_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [63:0] deq_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [1:0] deq_io_deq_bits_resp; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_bits_last; // @[Decoupled.scala 361:21]
  wire [29:0] deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  deq_metaReset; // @[Decoupled.scala 361:21]
  wire  q_b_deq_clock; // @[Decoupled.scala 361:21]
  wire  q_b_deq_reset; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] q_b_deq_io_enq_bits_id; // @[Decoupled.scala 361:21]
  wire [1:0] q_b_deq_io_enq_bits_resp; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_b_deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] q_b_deq_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [1:0] q_b_deq_io_deq_bits_resp; // @[Decoupled.scala 361:21]
  wire [29:0] q_b_deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  q_b_deq_metaReset; // @[Decoupled.scala 361:21]
  wire [15:0] _r_size1_T = {auto_in_ar_bits_len,8'hff}; // @[Cat.scala 31:58]
  wire [22:0] _GEN_0 = {{7'd0}, _r_size1_T}; // @[Bundles.scala 31:21]
  wire [22:0] _r_size1_T_1 = _GEN_0 << auto_in_ar_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] r_size1 = _r_size1_T_1[22:8]; // @[Bundles.scala 31:30]
  wire [15:0] _r_size_T = {r_size1, 1'h0}; // @[package.scala 232:35]
  wire [15:0] _r_size_T_1 = _r_size_T | 16'h1; // @[package.scala 232:40]
  wire [15:0] _r_size_T_2 = {1'h0,r_size1}; // @[Cat.scala 31:58]
  wire [15:0] _r_size_T_3 = ~_r_size_T_2; // @[package.scala 232:53]
  wire [15:0] _r_size_T_4 = _r_size_T_1 & _r_size_T_3; // @[package.scala 232:51]
  wire [7:0] r_size_hi = _r_size_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] r_size_lo = _r_size_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  _r_size_T_5 = |r_size_hi; // @[OneHot.scala 32:14]
  wire [7:0] _r_size_T_6 = r_size_hi | r_size_lo; // @[OneHot.scala 32:28]
  wire [3:0] r_size_hi_1 = _r_size_T_6[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] r_size_lo_1 = _r_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _r_size_T_7 = |r_size_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _r_size_T_8 = r_size_hi_1 | r_size_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] r_size_hi_2 = _r_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] r_size_lo_2 = _r_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _r_size_T_9 = |r_size_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _r_size_T_10 = r_size_hi_2 | r_size_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] r_size = {_r_size_T_5,_r_size_T_7,_r_size_T_9,_r_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  _r_ok_T_1 = r_size <= 4'hc; // @[Parameters.scala 92:42]
  wire [31:0] _r_ok_T_4 = auto_in_ar_bits_addr ^ 32'h3000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_5 = {1'b0,$signed(_r_ok_T_4)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_7 = $signed(_r_ok_T_5) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_8 = $signed(_r_ok_T_7) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _r_ok_T_9 = _r_ok_T_1 & _r_ok_T_8; // @[Parameters.scala 670:56]
  wire  _r_ok_T_11 = r_size <= 4'h6; // @[Parameters.scala 92:42]
  wire [32:0] _r_ok_T_15 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_17 = $signed(_r_ok_T_15) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_18 = $signed(_r_ok_T_17) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_19 = auto_in_ar_bits_addr ^ 32'h10000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_20 = {1'b0,$signed(_r_ok_T_19)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_22 = $signed(_r_ok_T_20) & -33'sh10000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_23 = $signed(_r_ok_T_22) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_24 = auto_in_ar_bits_addr ^ 32'h20000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_25 = {1'b0,$signed(_r_ok_T_24)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_27 = $signed(_r_ok_T_25) & -33'sh2000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_28 = $signed(_r_ok_T_27) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_29 = auto_in_ar_bits_addr ^ 32'h2000000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_30 = {1'b0,$signed(_r_ok_T_29)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_32 = $signed(_r_ok_T_30) & -33'sh10000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_33 = $signed(_r_ok_T_32) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_34 = auto_in_ar_bits_addr ^ 32'hc000000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_35 = {1'b0,$signed(_r_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_37 = $signed(_r_ok_T_35) & -33'sh4000000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_38 = $signed(_r_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_39 = auto_in_ar_bits_addr ^ 32'h64000000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_40 = {1'b0,$signed(_r_ok_T_39)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_42 = $signed(_r_ok_T_40) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_43 = $signed(_r_ok_T_42) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _r_ok_T_44 = auto_in_ar_bits_addr ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _r_ok_T_45 = {1'b0,$signed(_r_ok_T_44)}; // @[Parameters.scala 137:49]
  wire [32:0] _r_ok_T_47 = $signed(_r_ok_T_45) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _r_ok_T_48 = $signed(_r_ok_T_47) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _r_ok_T_54 = _r_ok_T_18 | _r_ok_T_23 | _r_ok_T_28 | _r_ok_T_33 | _r_ok_T_38 | _r_ok_T_43 | _r_ok_T_48; // @[Parameters.scala 671:42]
  wire  _r_ok_T_55 = _r_ok_T_11 & _r_ok_T_54; // @[Parameters.scala 670:56]
  wire  r_ok = _r_ok_T_9 | _r_ok_T_55; // @[Parameters.scala 672:30]
  wire [13:0] _GEN_114 = {{11'd0}, auto_in_ar_bits_addr[2:0]}; // @[ToTL.scala 90:59]
  wire [13:0] _r_addr_T_1 = 14'h3000 | _GEN_114; // @[ToTL.scala 90:59]
  wire [31:0] r_addr = r_ok ? auto_in_ar_bits_addr : {{18'd0}, _r_addr_T_1}; // @[ToTL.scala 90:23]
  reg [1:0] r_count_0; // @[ToTL.scala 91:28]
  reg [1:0] r_count_1; // @[ToTL.scala 91:28]
  reg [1:0] r_count_2; // @[ToTL.scala 91:28]
  reg [1:0] r_count_3; // @[ToTL.scala 91:28]
  reg [1:0] r_count_4; // @[ToTL.scala 91:28]
  reg [1:0] r_count_5; // @[ToTL.scala 91:28]
  reg [1:0] r_count_6; // @[ToTL.scala 91:28]
  reg [1:0] r_count_7; // @[ToTL.scala 91:28]
  reg [1:0] r_count_8; // @[ToTL.scala 91:28]
  reg [1:0] r_count_9; // @[ToTL.scala 91:28]
  reg [1:0] r_count_10; // @[ToTL.scala 91:28]
  reg [1:0] r_count_11; // @[ToTL.scala 91:28]
  reg [1:0] r_count_12; // @[ToTL.scala 91:28]
  reg [1:0] r_count_13; // @[ToTL.scala 91:28]
  reg [1:0] r_count_14; // @[ToTL.scala 91:28]
  reg [1:0] r_count_15; // @[ToTL.scala 91:28]
  wire [1:0] _GEN_1 = 4'h1 == auto_in_ar_bits_id ? r_count_1 : r_count_0; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_2 = 4'h2 == auto_in_ar_bits_id ? r_count_2 : _GEN_1; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_3 = 4'h3 == auto_in_ar_bits_id ? r_count_3 : _GEN_2; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_4 = 4'h4 == auto_in_ar_bits_id ? r_count_4 : _GEN_3; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_5 = 4'h5 == auto_in_ar_bits_id ? r_count_5 : _GEN_4; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_6 = 4'h6 == auto_in_ar_bits_id ? r_count_6 : _GEN_5; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_7 = 4'h7 == auto_in_ar_bits_id ? r_count_7 : _GEN_6; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_8 = 4'h8 == auto_in_ar_bits_id ? r_count_8 : _GEN_7; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_9 = 4'h9 == auto_in_ar_bits_id ? r_count_9 : _GEN_8; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_10 = 4'ha == auto_in_ar_bits_id ? r_count_10 : _GEN_9; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_11 = 4'hb == auto_in_ar_bits_id ? r_count_11 : _GEN_10; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_12 = 4'hc == auto_in_ar_bits_id ? r_count_12 : _GEN_11; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_13 = 4'hd == auto_in_ar_bits_id ? r_count_13 : _GEN_12; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_14 = 4'he == auto_in_ar_bits_id ? r_count_14 : _GEN_13; // @[ToTL.scala 95:{50,50}]
  wire [1:0] _GEN_15 = 4'hf == auto_in_ar_bits_id ? r_count_15 : _GEN_14; // @[ToTL.scala 95:{50,50}]
  wire [5:0] r_id = {auto_in_ar_bits_id,_GEN_15[0],1'h0}; // @[Cat.scala 31:58]
  wire [29:0] _T_2 = 30'h7fff << r_size; // @[package.scala 234:77]
  wire [14:0] _T_4 = ~_T_2[14:0]; // @[package.scala 234:46]
  wire  _T_8 = ~reset; // @[ToTL.scala 98:14]
  wire [1:0] a_mask_sizeOH_shiftAmount = r_size[1:0]; // @[OneHot.scala 63:49]
  wire [3:0] _a_mask_sizeOH_T_1 = 4'h1 << a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [2:0] a_mask_sizeOH = _a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _a_mask_T = r_size >= 4'h3; // @[Misc.scala 205:21]
  wire  a_mask_size = a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  a_mask_bit = r_addr[2]; // @[Misc.scala 209:26]
  wire  a_mask_nbit = ~a_mask_bit; // @[Misc.scala 210:20]
  wire  a_mask_acc = _a_mask_T | a_mask_size & a_mask_nbit; // @[Misc.scala 214:29]
  wire  a_mask_acc_1 = _a_mask_T | a_mask_size & a_mask_bit; // @[Misc.scala 214:29]
  wire  a_mask_size_1 = a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  a_mask_bit_1 = r_addr[1]; // @[Misc.scala 209:26]
  wire  a_mask_nbit_1 = ~a_mask_bit_1; // @[Misc.scala 210:20]
  wire  a_mask_eq_2 = a_mask_nbit & a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_2 = a_mask_acc | a_mask_size_1 & a_mask_eq_2; // @[Misc.scala 214:29]
  wire  a_mask_eq_3 = a_mask_nbit & a_mask_bit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_3 = a_mask_acc | a_mask_size_1 & a_mask_eq_3; // @[Misc.scala 214:29]
  wire  a_mask_eq_4 = a_mask_bit & a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_4 = a_mask_acc_1 | a_mask_size_1 & a_mask_eq_4; // @[Misc.scala 214:29]
  wire  a_mask_eq_5 = a_mask_bit & a_mask_bit_1; // @[Misc.scala 213:27]
  wire  a_mask_acc_5 = a_mask_acc_1 | a_mask_size_1 & a_mask_eq_5; // @[Misc.scala 214:29]
  wire  a_mask_size_2 = a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  a_mask_bit_2 = r_addr[0]; // @[Misc.scala 209:26]
  wire  a_mask_nbit_2 = ~a_mask_bit_2; // @[Misc.scala 210:20]
  wire  a_mask_eq_6 = a_mask_eq_2 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_6 = a_mask_acc_2 | a_mask_size_2 & a_mask_eq_6; // @[Misc.scala 214:29]
  wire  a_mask_eq_7 = a_mask_eq_2 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_7 = a_mask_acc_2 | a_mask_size_2 & a_mask_eq_7; // @[Misc.scala 214:29]
  wire  a_mask_eq_8 = a_mask_eq_3 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_8 = a_mask_acc_3 | a_mask_size_2 & a_mask_eq_8; // @[Misc.scala 214:29]
  wire  a_mask_eq_9 = a_mask_eq_3 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_9 = a_mask_acc_3 | a_mask_size_2 & a_mask_eq_9; // @[Misc.scala 214:29]
  wire  a_mask_eq_10 = a_mask_eq_4 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_10 = a_mask_acc_4 | a_mask_size_2 & a_mask_eq_10; // @[Misc.scala 214:29]
  wire  a_mask_eq_11 = a_mask_eq_4 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_11 = a_mask_acc_4 | a_mask_size_2 & a_mask_eq_11; // @[Misc.scala 214:29]
  wire  a_mask_eq_12 = a_mask_eq_5 & a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_12 = a_mask_acc_5 | a_mask_size_2 & a_mask_eq_12; // @[Misc.scala 214:29]
  wire  a_mask_eq_13 = a_mask_eq_5 & a_mask_bit_2; // @[Misc.scala 213:27]
  wire  a_mask_acc_13 = a_mask_acc_5 | a_mask_size_2 & a_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] a_mask = {a_mask_acc_13,a_mask_acc_12,a_mask_acc_11,a_mask_acc_10,a_mask_acc_9,a_mask_acc_8,a_mask_acc_7,
    a_mask_acc_6}; // @[Cat.scala 31:58]
  wire  r_out_bits_user_amba_prot_privileged = auto_in_ar_bits_prot[0]; // @[ToTL.scala 105:45]
  wire  r_out_bits_user_amba_prot_secure = ~auto_in_ar_bits_prot[1]; // @[ToTL.scala 106:29]
  wire  r_out_bits_user_amba_prot_fetch = auto_in_ar_bits_prot[2]; // @[ToTL.scala 107:45]
  wire  r_out_bits_user_amba_prot_bufferable = auto_in_ar_bits_cache[0]; // @[ToTL.scala 108:46]
  wire  r_out_bits_user_amba_prot_modifiable = auto_in_ar_bits_cache[1]; // @[ToTL.scala 109:46]
  wire  r_out_bits_user_amba_prot_readalloc = auto_in_ar_bits_cache[2]; // @[ToTL.scala 110:46]
  wire  r_out_bits_user_amba_prot_writealloc = auto_in_ar_bits_cache[3]; // @[ToTL.scala 111:46]
  wire [15:0] r_sel = 16'h1 << auto_in_ar_bits_id; // @[OneHot.scala 64:12]
  reg [7:0] beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = beatsLeft == 8'h0; // @[Arbiter.scala 88:28]
  wire  w_out_valid = auto_in_aw_valid & auto_in_w_valid; // @[ToTL.scala 135:34]
  wire [1:0] readys_valid = {w_out_valid,auto_in_ar_valid}; // @[Cat.scala 31:58]
  reg [1:0] readys_mask; // @[Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[Arbiter.scala 24:30]
  wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter = {_readys_filter_T_1,w_out_valid,auto_in_ar_valid}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_115 = {{1'd0}, readys_filter[3:1]}; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_115; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_116 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready = _GEN_116 | _readys_unready_T_4; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 26:18]
  wire  readys_0 = readys_readys[0]; // @[Arbiter.scala 95:86]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  out_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 123:31]
  wire  _T_26 = out_ready & auto_in_ar_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _r_count_0_T_1 = r_count_0 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_1_T_1 = r_count_1 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_2_T_1 = r_count_2 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_3_T_1 = r_count_3 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_4_T_1 = r_count_4 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_5_T_1 = r_count_5 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_6_T_1 = r_count_6 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_7_T_1 = r_count_7 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_8_T_1 = r_count_8 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_9_T_1 = r_count_9 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_10_T_1 = r_count_10 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_11_T_1 = r_count_11 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_12_T_1 = r_count_12 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_13_T_1 = r_count_13 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_14_T_1 = r_count_14 + 2'h1; // @[ToTL.scala 116:43]
  wire [1:0] _r_count_15_T_1 = r_count_15 + 2'h1; // @[ToTL.scala 116:43]
  wire [15:0] _w_size1_T = {auto_in_aw_bits_len,8'hff}; // @[Cat.scala 31:58]
  wire [22:0] _GEN_65 = {{7'd0}, _w_size1_T}; // @[Bundles.scala 31:21]
  wire [22:0] _w_size1_T_1 = _GEN_65 << auto_in_aw_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] w_size1 = _w_size1_T_1[22:8]; // @[Bundles.scala 31:30]
  wire [15:0] _w_size_T = {w_size1, 1'h0}; // @[package.scala 232:35]
  wire [15:0] _w_size_T_1 = _w_size_T | 16'h1; // @[package.scala 232:40]
  wire [15:0] _w_size_T_2 = {1'h0,w_size1}; // @[Cat.scala 31:58]
  wire [15:0] _w_size_T_3 = ~_w_size_T_2; // @[package.scala 232:53]
  wire [15:0] _w_size_T_4 = _w_size_T_1 & _w_size_T_3; // @[package.scala 232:51]
  wire [7:0] w_size_hi = _w_size_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] w_size_lo = _w_size_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  _w_size_T_5 = |w_size_hi; // @[OneHot.scala 32:14]
  wire [7:0] _w_size_T_6 = w_size_hi | w_size_lo; // @[OneHot.scala 32:28]
  wire [3:0] w_size_hi_1 = _w_size_T_6[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] w_size_lo_1 = _w_size_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _w_size_T_7 = |w_size_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _w_size_T_8 = w_size_hi_1 | w_size_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] w_size_hi_2 = _w_size_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] w_size_lo_2 = _w_size_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _w_size_T_9 = |w_size_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _w_size_T_10 = w_size_hi_2 | w_size_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] w_size = {_w_size_T_5,_w_size_T_7,_w_size_T_9,_w_size_T_10[1]}; // @[Cat.scala 31:58]
  wire  _w_ok_T_1 = w_size <= 4'hc; // @[Parameters.scala 92:42]
  wire [31:0] _w_ok_T_4 = auto_in_aw_bits_addr ^ 32'h3000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_5 = {1'b0,$signed(_w_ok_T_4)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_7 = $signed(_w_ok_T_5) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_8 = $signed(_w_ok_T_7) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _w_ok_T_9 = _w_ok_T_1 & _w_ok_T_8; // @[Parameters.scala 670:56]
  wire  _w_ok_T_11 = w_size <= 4'h6; // @[Parameters.scala 92:42]
  wire [32:0] _w_ok_T_15 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_17 = $signed(_w_ok_T_15) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_18 = $signed(_w_ok_T_17) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _w_ok_T_19 = auto_in_aw_bits_addr ^ 32'h2000000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_20 = {1'b0,$signed(_w_ok_T_19)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_22 = $signed(_w_ok_T_20) & -33'sh10000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_23 = $signed(_w_ok_T_22) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _w_ok_T_24 = auto_in_aw_bits_addr ^ 32'hc000000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_25 = {1'b0,$signed(_w_ok_T_24)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_27 = $signed(_w_ok_T_25) & -33'sh4000000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_28 = $signed(_w_ok_T_27) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _w_ok_T_29 = auto_in_aw_bits_addr ^ 32'h64000000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_30 = {1'b0,$signed(_w_ok_T_29)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_32 = $signed(_w_ok_T_30) & -33'sh1000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_33 = $signed(_w_ok_T_32) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _w_ok_T_34 = auto_in_aw_bits_addr ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _w_ok_T_35 = {1'b0,$signed(_w_ok_T_34)}; // @[Parameters.scala 137:49]
  wire [32:0] _w_ok_T_37 = $signed(_w_ok_T_35) & -33'sh80000000; // @[Parameters.scala 137:52]
  wire  _w_ok_T_38 = $signed(_w_ok_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _w_ok_T_42 = _w_ok_T_18 | _w_ok_T_23 | _w_ok_T_28 | _w_ok_T_33 | _w_ok_T_38; // @[Parameters.scala 671:42]
  wire  _w_ok_T_43 = _w_ok_T_11 & _w_ok_T_42; // @[Parameters.scala 670:56]
  wire  w_ok = _w_ok_T_9 | _w_ok_T_43; // @[Parameters.scala 672:30]
  wire [13:0] _GEN_117 = {{11'd0}, auto_in_aw_bits_addr[2:0]}; // @[ToTL.scala 123:59]
  wire [13:0] _w_addr_T_1 = 14'h3000 | _GEN_117; // @[ToTL.scala 123:59]
  wire [31:0] w_addr = w_ok ? auto_in_aw_bits_addr : {{18'd0}, _w_addr_T_1}; // @[ToTL.scala 123:23]
  reg [1:0] w_count_0; // @[ToTL.scala 124:28]
  reg [1:0] w_count_1; // @[ToTL.scala 124:28]
  reg [1:0] w_count_2; // @[ToTL.scala 124:28]
  reg [1:0] w_count_3; // @[ToTL.scala 124:28]
  reg [1:0] w_count_4; // @[ToTL.scala 124:28]
  reg [1:0] w_count_5; // @[ToTL.scala 124:28]
  reg [1:0] w_count_6; // @[ToTL.scala 124:28]
  reg [1:0] w_count_7; // @[ToTL.scala 124:28]
  reg [1:0] w_count_8; // @[ToTL.scala 124:28]
  reg [1:0] w_count_9; // @[ToTL.scala 124:28]
  reg [1:0] w_count_10; // @[ToTL.scala 124:28]
  reg [1:0] w_count_11; // @[ToTL.scala 124:28]
  reg [1:0] w_count_12; // @[ToTL.scala 124:28]
  reg [1:0] w_count_13; // @[ToTL.scala 124:28]
  reg [1:0] w_count_14; // @[ToTL.scala 124:28]
  reg [1:0] w_count_15; // @[ToTL.scala 124:28]
  wire [1:0] _GEN_33 = 4'h1 == auto_in_aw_bits_id ? w_count_1 : w_count_0; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_34 = 4'h2 == auto_in_aw_bits_id ? w_count_2 : _GEN_33; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_35 = 4'h3 == auto_in_aw_bits_id ? w_count_3 : _GEN_34; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_36 = 4'h4 == auto_in_aw_bits_id ? w_count_4 : _GEN_35; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_37 = 4'h5 == auto_in_aw_bits_id ? w_count_5 : _GEN_36; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_38 = 4'h6 == auto_in_aw_bits_id ? w_count_6 : _GEN_37; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_39 = 4'h7 == auto_in_aw_bits_id ? w_count_7 : _GEN_38; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_40 = 4'h8 == auto_in_aw_bits_id ? w_count_8 : _GEN_39; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_41 = 4'h9 == auto_in_aw_bits_id ? w_count_9 : _GEN_40; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_42 = 4'ha == auto_in_aw_bits_id ? w_count_10 : _GEN_41; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_43 = 4'hb == auto_in_aw_bits_id ? w_count_11 : _GEN_42; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_44 = 4'hc == auto_in_aw_bits_id ? w_count_12 : _GEN_43; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_45 = 4'hd == auto_in_aw_bits_id ? w_count_13 : _GEN_44; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_46 = 4'he == auto_in_aw_bits_id ? w_count_14 : _GEN_45; // @[ToTL.scala 128:{50,50}]
  wire [1:0] _GEN_47 = 4'hf == auto_in_aw_bits_id ? w_count_15 : _GEN_46; // @[ToTL.scala 128:{50,50}]
  wire [5:0] w_id = {auto_in_aw_bits_id,_GEN_47[0],1'h1}; // @[Cat.scala 31:58]
  wire  _T_58 = ~auto_in_aw_valid; // @[ToTL.scala 131:15]
  wire [29:0] _T_60 = 30'h7fff << w_size; // @[package.scala 234:77]
  wire [14:0] _T_62 = ~_T_60[14:0]; // @[package.scala 234:46]
  wire  readys_1 = readys_readys[1]; // @[Arbiter.scala 95:86]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire  out_1_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 123:31]
  wire  bundleIn_0_aw_ready = out_1_ready & auto_in_w_valid & auto_in_w_bits_last; // @[ToTL.scala 133:48]
  wire  w_out_bits_user_amba_prot_privileged = auto_in_aw_bits_prot[0]; // @[ToTL.scala 141:45]
  wire  w_out_bits_user_amba_prot_secure = ~auto_in_aw_bits_prot[1]; // @[ToTL.scala 142:29]
  wire  w_out_bits_user_amba_prot_fetch = auto_in_aw_bits_prot[2]; // @[ToTL.scala 143:45]
  wire  w_out_bits_user_amba_prot_bufferable = auto_in_aw_bits_cache[0]; // @[ToTL.scala 144:46]
  wire  w_out_bits_user_amba_prot_modifiable = auto_in_aw_bits_cache[1]; // @[ToTL.scala 145:46]
  wire  w_out_bits_user_amba_prot_readalloc = auto_in_aw_bits_cache[2]; // @[ToTL.scala 146:46]
  wire  w_out_bits_user_amba_prot_writealloc = auto_in_aw_bits_cache[3]; // @[ToTL.scala 147:46]
  wire [15:0] w_sel = 16'h1 << auto_in_aw_bits_id; // @[OneHot.scala 64:12]
  wire  _T_92 = bundleIn_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _w_count_0_T_1 = w_count_0 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_1_T_1 = w_count_1 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_2_T_1 = w_count_2 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_3_T_1 = w_count_3 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_4_T_1 = w_count_4 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_5_T_1 = w_count_5 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_6_T_1 = w_count_6 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_7_T_1 = w_count_7 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_8_T_1 = w_count_8 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_9_T_1 = w_count_9 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_10_T_1 = w_count_10 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_11_T_1 = w_count_11 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_12_T_1 = w_count_12 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_13_T_1 = w_count_13 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_14_T_1 = w_count_14 + 2'h1; // @[ToTL.scala 152:43]
  wire [1:0] _w_count_15_T_1 = w_count_15 + 2'h1; // @[ToTL.scala 152:43]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 89:24]
  wire [1:0] _readys_mask_T = readys_readys & readys_valid; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[package.scala 244:43]
  wire  earlyWinner_0 = readys_0 & auto_in_ar_valid; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1 = readys_1 & w_out_valid; // @[Arbiter.scala 97:79]
  wire  _T_134 = auto_in_ar_valid | w_out_valid; // @[Arbiter.scala 107:36]
  wire  _T_135 = ~(auto_in_ar_valid | w_out_valid); // @[Arbiter.scala 107:15]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & auto_in_ar_valid | state_1 & w_out_valid; // @[Mux.scala 27:73]
  wire  sink_ACancel_earlyValid = idle ? _T_134 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire [7:0] _GEN_118 = {{7'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  wire [7:0] _beatsLeft_T_4 = beatsLeft - _GEN_118; // @[Arbiter.scala 113:52]
  wire [7:0] _T_154 = muxStateEarly_0 ? a_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _T_155 = muxStateEarly_1 ? auto_in_w_bits_strb : 8'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_178 = muxStateEarly_0 ? r_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_179 = muxStateEarly_1 ? w_addr : 32'h0; // @[Mux.scala 27:73]
  wire [5:0] _T_181 = muxStateEarly_0 ? r_id : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _T_182 = muxStateEarly_1 ? w_id : 6'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_184 = muxStateEarly_0 ? r_size : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_185 = muxStateEarly_1 ? w_size : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_190 = muxStateEarly_0 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_191 = muxStateEarly_1 ? 3'h1 : 3'h0; // @[Mux.scala 27:73]
  wire  d_hasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  ok_r_ready = deq_io_enq_ready; // @[ToTL.scala 158:23 Decoupled.scala 365:17]
  wire  ok_b_ready = q_b_deq_io_enq_ready; // @[ToTL.scala 157:23 Decoupled.scala 365:17]
  wire  bundleOut_0_d_ready = d_hasData ? ok_r_ready : ok_b_ready; // @[ToTL.scala 164:25]
  wire  _d_last_T = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 50:35]
  wire [26:0] _d_last_beats1_decode_T_1 = 27'hfff << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [11:0] _d_last_beats1_decode_T_3 = ~_d_last_beats1_decode_T_1[11:0]; // @[package.scala 234:46]
  wire [8:0] d_last_beats1_decode = _d_last_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59]
  wire [8:0] d_last_beats1 = d_hasData ? d_last_beats1_decode : 9'h0; // @[Edges.scala 220:14]
  reg [8:0] d_last_counter; // @[Edges.scala 228:27]
  wire [8:0] d_last_counter1 = d_last_counter - 9'h1; // @[Edges.scala 229:28]
  wire  d_last_first = d_last_counter == 9'h0; // @[Edges.scala 230:25]
  reg [1:0] b_count_0; // @[ToTL.scala 186:28]
  reg [1:0] b_count_1; // @[ToTL.scala 186:28]
  reg [1:0] b_count_2; // @[ToTL.scala 186:28]
  reg [1:0] b_count_3; // @[ToTL.scala 186:28]
  reg [1:0] b_count_4; // @[ToTL.scala 186:28]
  reg [1:0] b_count_5; // @[ToTL.scala 186:28]
  reg [1:0] b_count_6; // @[ToTL.scala 186:28]
  reg [1:0] b_count_7; // @[ToTL.scala 186:28]
  reg [1:0] b_count_8; // @[ToTL.scala 186:28]
  reg [1:0] b_count_9; // @[ToTL.scala 186:28]
  reg [1:0] b_count_10; // @[ToTL.scala 186:28]
  reg [1:0] b_count_11; // @[ToTL.scala 186:28]
  reg [1:0] b_count_12; // @[ToTL.scala 186:28]
  reg [1:0] b_count_13; // @[ToTL.scala 186:28]
  reg [1:0] b_count_14; // @[ToTL.scala 186:28]
  reg [1:0] b_count_15; // @[ToTL.scala 186:28]
  wire [3:0] q_b_bits_id = q_b_deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  wire [1:0] _GEN_67 = 4'h1 == q_b_bits_id ? b_count_1 : b_count_0; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_68 = 4'h2 == q_b_bits_id ? b_count_2 : _GEN_67; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_69 = 4'h3 == q_b_bits_id ? b_count_3 : _GEN_68; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_70 = 4'h4 == q_b_bits_id ? b_count_4 : _GEN_69; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_71 = 4'h5 == q_b_bits_id ? b_count_5 : _GEN_70; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_72 = 4'h6 == q_b_bits_id ? b_count_6 : _GEN_71; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_73 = 4'h7 == q_b_bits_id ? b_count_7 : _GEN_72; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_74 = 4'h8 == q_b_bits_id ? b_count_8 : _GEN_73; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_75 = 4'h9 == q_b_bits_id ? b_count_9 : _GEN_74; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_76 = 4'ha == q_b_bits_id ? b_count_10 : _GEN_75; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_77 = 4'hb == q_b_bits_id ? b_count_11 : _GEN_76; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_78 = 4'hc == q_b_bits_id ? b_count_12 : _GEN_77; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_79 = 4'hd == q_b_bits_id ? b_count_13 : _GEN_78; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_80 = 4'he == q_b_bits_id ? b_count_14 : _GEN_79; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_81 = 4'hf == q_b_bits_id ? b_count_15 : _GEN_80; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_83 = 4'h1 == q_b_bits_id ? w_count_1 : w_count_0; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_84 = 4'h2 == q_b_bits_id ? w_count_2 : _GEN_83; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_85 = 4'h3 == q_b_bits_id ? w_count_3 : _GEN_84; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_86 = 4'h4 == q_b_bits_id ? w_count_4 : _GEN_85; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_87 = 4'h5 == q_b_bits_id ? w_count_5 : _GEN_86; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_88 = 4'h6 == q_b_bits_id ? w_count_6 : _GEN_87; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_89 = 4'h7 == q_b_bits_id ? w_count_7 : _GEN_88; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_90 = 4'h8 == q_b_bits_id ? w_count_8 : _GEN_89; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_91 = 4'h9 == q_b_bits_id ? w_count_9 : _GEN_90; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_92 = 4'ha == q_b_bits_id ? w_count_10 : _GEN_91; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_93 = 4'hb == q_b_bits_id ? w_count_11 : _GEN_92; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_94 = 4'hc == q_b_bits_id ? w_count_12 : _GEN_93; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_95 = 4'hd == q_b_bits_id ? w_count_13 : _GEN_94; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_96 = 4'he == q_b_bits_id ? w_count_14 : _GEN_95; // @[ToTL.scala 187:{43,43}]
  wire [1:0] _GEN_97 = 4'hf == q_b_bits_id ? w_count_15 : _GEN_96; // @[ToTL.scala 187:{43,43}]
  wire  b_allow = _GEN_81 != _GEN_97; // @[ToTL.scala 187:43]
  wire [15:0] b_sel = 16'h1 << q_b_bits_id; // @[OneHot.scala 64:12]
  wire  q_b_valid = q_b_deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  wire  bundleIn_0_b_valid = q_b_valid & b_allow; // @[ToTL.scala 195:31]
  wire  _T_209 = auto_in_b_ready & bundleIn_0_b_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _b_count_0_T_1 = b_count_0 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_1_T_1 = b_count_1 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_2_T_1 = b_count_2 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_3_T_1 = b_count_3 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_4_T_1 = b_count_4 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_5_T_1 = b_count_5 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_6_T_1 = b_count_6 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_7_T_1 = b_count_7 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_8_T_1 = b_count_8 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_9_T_1 = b_count_9 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_10_T_1 = b_count_10 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_11_T_1 = b_count_11 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_12_T_1 = b_count_12 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_13_T_1 = b_count_13 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_14_T_1 = b_count_14 + 2'h1; // @[ToTL.scala 191:42]
  wire [1:0] _b_count_15_T_1 = b_count_15 + 2'h1; // @[ToTL.scala 191:42]
  reg [6:0] AXI4ToTL_1_covState; // @[Register tracking AXI4ToTL_1 state]
  reg  AXI4ToTL_1_covMap [0:127]; // @[Coverage map for AXI4ToTL_1]
  wire  AXI4ToTL_1_covMap_read_en; // @[Coverage map for AXI4ToTL_1]
  wire [6:0] AXI4ToTL_1_covMap_read_addr; // @[Coverage map for AXI4ToTL_1]
  wire  AXI4ToTL_1_covMap_read_data; // @[Coverage map for AXI4ToTL_1]
  wire  AXI4ToTL_1_covMap_write_data; // @[Coverage map for AXI4ToTL_1]
  wire [6:0] AXI4ToTL_1_covMap_write_addr; // @[Coverage map for AXI4ToTL_1]
  wire  AXI4ToTL_1_covMap_write_mask; // @[Coverage map for AXI4ToTL_1]
  wire  AXI4ToTL_1_covMap_write_en; // @[Coverage map for AXI4ToTL_1]
  reg [29:0] AXI4ToTL_1_covSum; // @[Sum of coverage map]
  wire [1:0] readys_mask_shl;
  wire [6:0] readys_mask_pad;
  wire [3:0] w_count_4_shl;
  wire [6:0] w_count_4_pad;
  wire [3:0] w_count_14_shl;
  wire [6:0] w_count_14_pad;
  wire [6:0] b_count_5_shl;
  wire [6:0] b_count_5_pad;
  wire [6:0] b_count_3_shl;
  wire [6:0] b_count_3_pad;
  wire [3:0] w_count_7_shl;
  wire [6:0] w_count_7_pad;
  wire [3:0] w_count_3_shl;
  wire [6:0] w_count_3_pad;
  wire [6:0] b_count_10_shl;
  wire [6:0] b_count_10_pad;
  wire [3:0] w_count_1_shl;
  wire [6:0] w_count_1_pad;
  wire [3:0] w_count_2_shl;
  wire [6:0] w_count_2_pad;
  wire [6:0] b_count_11_shl;
  wire [6:0] b_count_11_pad;
  wire [6:0] b_count_7_shl;
  wire [6:0] b_count_7_pad;
  wire [6:0] b_count_8_shl;
  wire [6:0] b_count_8_pad;
  wire [6:0] b_count_13_shl;
  wire [6:0] b_count_13_pad;
  wire [3:0] w_count_12_shl;
  wire [6:0] w_count_12_pad;
  wire [6:0] b_count_6_shl;
  wire [6:0] b_count_6_pad;
  wire [3:0] w_count_10_shl;
  wire [6:0] w_count_10_pad;
  wire [3:0] w_count_9_shl;
  wire [6:0] w_count_9_pad;
  wire [3:0] w_count_6_shl;
  wire [6:0] w_count_6_pad;
  wire [6:0] b_count_4_shl;
  wire [6:0] b_count_4_pad;
  wire [6:0] b_count_14_shl;
  wire [6:0] b_count_14_pad;
  wire [6:0] b_count_2_shl;
  wire [6:0] b_count_2_pad;
  wire [6:0] b_count_1_shl;
  wire [6:0] b_count_1_pad;
  wire [3:0] w_count_8_shl;
  wire [6:0] w_count_8_pad;
  wire [6:0] b_count_0_shl;
  wire [6:0] b_count_0_pad;
  wire [4:0] state_1_shl;
  wire [6:0] state_1_pad;
  wire [4:0] state_0_shl;
  wire [6:0] state_0_pad;
  wire [3:0] w_count_15_shl;
  wire [6:0] w_count_15_pad;
  wire [6:0] b_count_12_shl;
  wire [6:0] b_count_12_pad;
  wire [3:0] w_count_11_shl;
  wire [6:0] w_count_11_pad;
  wire [6:0] b_count_9_shl;
  wire [6:0] b_count_9_pad;
  wire [3:0] w_count_13_shl;
  wire [6:0] w_count_13_pad;
  wire [3:0] w_count_5_shl;
  wire [6:0] w_count_5_pad;
  wire [6:0] b_count_15_shl;
  wire [6:0] b_count_15_pad;
  wire [3:0] w_count_0_shl;
  wire [6:0] w_count_0_pad;
  wire [6:0] AXI4ToTL_1_xor15;
  wire [6:0] AXI4ToTL_1_xor16;
  wire [6:0] AXI4ToTL_1_xor7;
  wire [6:0] AXI4ToTL_1_xor17;
  wire [6:0] AXI4ToTL_1_xor18;
  wire [6:0] AXI4ToTL_1_xor8;
  wire [6:0] AXI4ToTL_1_xor3;
  wire [6:0] AXI4ToTL_1_xor19;
  wire [6:0] AXI4ToTL_1_xor20;
  wire [6:0] AXI4ToTL_1_xor9;
  wire [6:0] AXI4ToTL_1_xor21;
  wire [6:0] AXI4ToTL_1_xor46;
  wire [6:0] AXI4ToTL_1_xor22;
  wire [6:0] AXI4ToTL_1_xor10;
  wire [6:0] AXI4ToTL_1_xor4;
  wire [6:0] AXI4ToTL_1_xor1;
  wire [6:0] AXI4ToTL_1_xor23;
  wire [6:0] AXI4ToTL_1_xor24;
  wire [6:0] AXI4ToTL_1_xor11;
  wire [6:0] AXI4ToTL_1_xor25;
  wire [6:0] AXI4ToTL_1_xor54;
  wire [6:0] AXI4ToTL_1_xor26;
  wire [6:0] AXI4ToTL_1_xor12;
  wire [6:0] AXI4ToTL_1_xor5;
  wire [6:0] AXI4ToTL_1_xor27;
  wire [6:0] AXI4ToTL_1_xor28;
  wire [6:0] AXI4ToTL_1_xor13;
  wire [6:0] AXI4ToTL_1_xor29;
  wire [6:0] AXI4ToTL_1_xor62;
  wire [6:0] AXI4ToTL_1_xor30;
  wire [6:0] AXI4ToTL_1_xor14;
  wire [6:0] AXI4ToTL_1_xor6;
  wire [6:0] AXI4ToTL_1_xor2;
  wire [6:0] AXI4ToTL_1_xor0;
  wire [29:0] deq_sum;
  wire [29:0] q_b_deq_sum;
  Queue_26 deq ( // @[Decoupled.scala 361:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_id(deq_io_enq_bits_id),
    .io_enq_bits_data(deq_io_enq_bits_data),
    .io_enq_bits_resp(deq_io_enq_bits_resp),
    .io_enq_bits_last(deq_io_enq_bits_last),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_id(deq_io_deq_bits_id),
    .io_deq_bits_data(deq_io_deq_bits_data),
    .io_deq_bits_resp(deq_io_deq_bits_resp),
    .io_deq_bits_last(deq_io_deq_bits_last),
    .io_covSum(deq_io_covSum),
    .metaReset(deq_metaReset)
  );
  Queue_27 q_b_deq ( // @[Decoupled.scala 361:21]
    .clock(q_b_deq_clock),
    .reset(q_b_deq_reset),
    .io_enq_ready(q_b_deq_io_enq_ready),
    .io_enq_valid(q_b_deq_io_enq_valid),
    .io_enq_bits_id(q_b_deq_io_enq_bits_id),
    .io_enq_bits_resp(q_b_deq_io_enq_bits_resp),
    .io_deq_ready(q_b_deq_io_deq_ready),
    .io_deq_valid(q_b_deq_io_deq_valid),
    .io_deq_bits_id(q_b_deq_io_deq_bits_id),
    .io_deq_bits_resp(q_b_deq_io_deq_bits_resp),
    .io_covSum(q_b_deq_io_covSum),
    .metaReset(q_b_deq_metaReset)
  );
  assign auto_in_aw_ready = out_1_ready & auto_in_w_valid & auto_in_w_bits_last; // @[ToTL.scala 133:48]
  assign auto_in_w_ready = out_1_ready & auto_in_aw_valid; // @[ToTL.scala 134:34]
  assign auto_in_b_valid = q_b_valid & b_allow; // @[ToTL.scala 195:31]
  assign auto_in_b_bits_id = q_b_deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_b_bits_resp = q_b_deq_io_deq_bits_resp; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_ar_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 123:31]
  assign auto_in_r_valid = deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  assign auto_in_r_bits_id = deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_r_bits_data = deq_io_deq_bits_data; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_r_bits_resp = deq_io_deq_bits_resp; // @[Decoupled.scala 401:19 402:14]
  assign auto_in_r_bits_last = deq_io_deq_bits_last; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_a_valid = idle ? _T_134 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign auto_out_a_bits_opcode = _T_190 | _T_191; // @[Mux.scala 27:73]
  assign auto_out_a_bits_size = _T_184 | _T_185; // @[Mux.scala 27:73]
  assign auto_out_a_bits_source = _T_181 | _T_182; // @[Mux.scala 27:73]
  assign auto_out_a_bits_address = _T_178 | _T_179; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_bufferable = muxStateEarly_0 & r_out_bits_user_amba_prot_bufferable |
    muxStateEarly_1 & w_out_bits_user_amba_prot_bufferable; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_modifiable = muxStateEarly_0 & r_out_bits_user_amba_prot_modifiable |
    muxStateEarly_1 & w_out_bits_user_amba_prot_modifiable; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_readalloc = muxStateEarly_0 & r_out_bits_user_amba_prot_readalloc |
    muxStateEarly_1 & w_out_bits_user_amba_prot_readalloc; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_writealloc = muxStateEarly_0 & r_out_bits_user_amba_prot_writealloc |
    muxStateEarly_1 & w_out_bits_user_amba_prot_writealloc; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_privileged = muxStateEarly_0 & r_out_bits_user_amba_prot_privileged |
    muxStateEarly_1 & w_out_bits_user_amba_prot_privileged; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_secure = muxStateEarly_0 & r_out_bits_user_amba_prot_secure | muxStateEarly_1 &
    w_out_bits_user_amba_prot_secure; // @[Mux.scala 27:73]
  assign auto_out_a_bits_user_amba_prot_fetch = muxStateEarly_0 & r_out_bits_user_amba_prot_fetch | muxStateEarly_1 &
    w_out_bits_user_amba_prot_fetch; // @[Mux.scala 27:73]
  assign auto_out_a_bits_mask = _T_154 | _T_155; // @[Mux.scala 27:73]
  assign auto_out_a_bits_data = muxStateEarly_1 ? auto_in_w_bits_data : 64'h0; // @[Mux.scala 27:73]
  assign auto_out_d_ready = d_hasData ? ok_r_ready : ok_b_ready; // @[ToTL.scala 164:25]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = auto_out_d_valid & d_hasData; // @[ToTL.scala 165:33]
  assign deq_io_enq_bits_id = auto_out_d_bits_source[5:2]; // @[ToTL.scala 168:43]
  assign deq_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign deq_io_enq_bits_resp = auto_out_d_bits_denied | auto_out_d_bits_corrupt ? 2'h2 : 2'h0; // @[ToTL.scala 160:23]
  assign deq_io_enq_bits_last = d_last_counter == 9'h1 | d_last_beats1 == 9'h0; // @[Edges.scala 231:37]
  assign deq_io_deq_ready = auto_in_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign q_b_deq_clock = clock;
  assign q_b_deq_reset = reset;
  assign q_b_deq_io_enq_valid = auto_out_d_valid & ~d_hasData; // @[ToTL.scala 166:33]
  assign q_b_deq_io_enq_bits_id = auto_out_d_bits_source[5:2]; // @[ToTL.scala 177:43]
  assign q_b_deq_io_enq_bits_resp = auto_out_d_bits_denied | auto_out_d_bits_corrupt ? 2'h2 : 2'h0; // @[ToTL.scala 160:23]
  assign q_b_deq_io_deq_ready = auto_in_b_ready & b_allow; // @[ToTL.scala 196:31]
  assign AXI4ToTL_1_covMap_read_en = 1'h1;
  assign AXI4ToTL_1_covMap_read_addr = AXI4ToTL_1_covState;
  assign AXI4ToTL_1_covMap_read_data = AXI4ToTL_1_covMap[AXI4ToTL_1_covMap_read_addr]; // @[Coverage map for AXI4ToTL_1]
  assign AXI4ToTL_1_covMap_write_data = 1'h1;
  assign AXI4ToTL_1_covMap_write_addr = AXI4ToTL_1_covState;
  assign AXI4ToTL_1_covMap_write_mask = 1'h1;
  assign AXI4ToTL_1_covMap_write_en = ~metaReset;
  assign readys_mask_shl = readys_mask;
  assign readys_mask_pad = {5'h0,readys_mask_shl};
  assign w_count_4_shl = {w_count_4, 2'h0};
  assign w_count_4_pad = {3'h0,w_count_4_shl};
  assign w_count_14_shl = {w_count_14, 2'h0};
  assign w_count_14_pad = {3'h0,w_count_14_shl};
  assign b_count_5_shl = {b_count_5, 5'h0};
  assign b_count_5_pad = b_count_5_shl;
  assign b_count_3_shl = {b_count_3, 5'h0};
  assign b_count_3_pad = b_count_3_shl;
  assign w_count_7_shl = {w_count_7, 2'h0};
  assign w_count_7_pad = {3'h0,w_count_7_shl};
  assign w_count_3_shl = {w_count_3, 2'h0};
  assign w_count_3_pad = {3'h0,w_count_3_shl};
  assign b_count_10_shl = {b_count_10, 5'h0};
  assign b_count_10_pad = b_count_10_shl;
  assign w_count_1_shl = {w_count_1, 2'h0};
  assign w_count_1_pad = {3'h0,w_count_1_shl};
  assign w_count_2_shl = {w_count_2, 2'h0};
  assign w_count_2_pad = {3'h0,w_count_2_shl};
  assign b_count_11_shl = {b_count_11, 5'h0};
  assign b_count_11_pad = b_count_11_shl;
  assign b_count_7_shl = {b_count_7, 5'h0};
  assign b_count_7_pad = b_count_7_shl;
  assign b_count_8_shl = {b_count_8, 5'h0};
  assign b_count_8_pad = b_count_8_shl;
  assign b_count_13_shl = {b_count_13, 5'h0};
  assign b_count_13_pad = b_count_13_shl;
  assign w_count_12_shl = {w_count_12, 2'h0};
  assign w_count_12_pad = {3'h0,w_count_12_shl};
  assign b_count_6_shl = {b_count_6, 5'h0};
  assign b_count_6_pad = b_count_6_shl;
  assign w_count_10_shl = {w_count_10, 2'h0};
  assign w_count_10_pad = {3'h0,w_count_10_shl};
  assign w_count_9_shl = {w_count_9, 2'h0};
  assign w_count_9_pad = {3'h0,w_count_9_shl};
  assign w_count_6_shl = {w_count_6, 2'h0};
  assign w_count_6_pad = {3'h0,w_count_6_shl};
  assign b_count_4_shl = {b_count_4, 5'h0};
  assign b_count_4_pad = b_count_4_shl;
  assign b_count_14_shl = {b_count_14, 5'h0};
  assign b_count_14_pad = b_count_14_shl;
  assign b_count_2_shl = {b_count_2, 5'h0};
  assign b_count_2_pad = b_count_2_shl;
  assign b_count_1_shl = {b_count_1, 5'h0};
  assign b_count_1_pad = b_count_1_shl;
  assign w_count_8_shl = {w_count_8, 2'h0};
  assign w_count_8_pad = {3'h0,w_count_8_shl};
  assign b_count_0_shl = {b_count_0, 5'h0};
  assign b_count_0_pad = b_count_0_shl;
  assign state_1_shl = {state_1, 4'h0};
  assign state_1_pad = {2'h0,state_1_shl};
  assign state_0_shl = {state_0, 4'h0};
  assign state_0_pad = {2'h0,state_0_shl};
  assign w_count_15_shl = {w_count_15, 2'h0};
  assign w_count_15_pad = {3'h0,w_count_15_shl};
  assign b_count_12_shl = {b_count_12, 5'h0};
  assign b_count_12_pad = b_count_12_shl;
  assign w_count_11_shl = {w_count_11, 2'h0};
  assign w_count_11_pad = {3'h0,w_count_11_shl};
  assign b_count_9_shl = {b_count_9, 5'h0};
  assign b_count_9_pad = b_count_9_shl;
  assign w_count_13_shl = {w_count_13, 2'h0};
  assign w_count_13_pad = {3'h0,w_count_13_shl};
  assign w_count_5_shl = {w_count_5, 2'h0};
  assign w_count_5_pad = {3'h0,w_count_5_shl};
  assign b_count_15_shl = {b_count_15, 5'h0};
  assign b_count_15_pad = b_count_15_shl;
  assign w_count_0_shl = {w_count_0, 2'h0};
  assign w_count_0_pad = {3'h0,w_count_0_shl};
  assign AXI4ToTL_1_xor15 = readys_mask_pad ^ w_count_4_pad;
  assign AXI4ToTL_1_xor16 = w_count_14_pad ^ b_count_5_pad;
  assign AXI4ToTL_1_xor7 = AXI4ToTL_1_xor15 ^ AXI4ToTL_1_xor16;
  assign AXI4ToTL_1_xor17 = b_count_3_pad ^ w_count_7_pad;
  assign AXI4ToTL_1_xor18 = w_count_3_pad ^ b_count_10_pad;
  assign AXI4ToTL_1_xor8 = AXI4ToTL_1_xor17 ^ AXI4ToTL_1_xor18;
  assign AXI4ToTL_1_xor3 = AXI4ToTL_1_xor7 ^ AXI4ToTL_1_xor8;
  assign AXI4ToTL_1_xor19 = w_count_1_pad ^ w_count_2_pad;
  assign AXI4ToTL_1_xor20 = b_count_11_pad ^ b_count_7_pad;
  assign AXI4ToTL_1_xor9 = AXI4ToTL_1_xor19 ^ AXI4ToTL_1_xor20;
  assign AXI4ToTL_1_xor21 = b_count_8_pad ^ b_count_13_pad;
  assign AXI4ToTL_1_xor46 = b_count_6_pad ^ w_count_10_pad;
  assign AXI4ToTL_1_xor22 = w_count_12_pad ^ AXI4ToTL_1_xor46;
  assign AXI4ToTL_1_xor10 = AXI4ToTL_1_xor21 ^ AXI4ToTL_1_xor22;
  assign AXI4ToTL_1_xor4 = AXI4ToTL_1_xor9 ^ AXI4ToTL_1_xor10;
  assign AXI4ToTL_1_xor1 = AXI4ToTL_1_xor3 ^ AXI4ToTL_1_xor4;
  assign AXI4ToTL_1_xor23 = w_count_9_pad ^ w_count_6_pad;
  assign AXI4ToTL_1_xor24 = b_count_4_pad ^ b_count_14_pad;
  assign AXI4ToTL_1_xor11 = AXI4ToTL_1_xor23 ^ AXI4ToTL_1_xor24;
  assign AXI4ToTL_1_xor25 = b_count_2_pad ^ b_count_1_pad;
  assign AXI4ToTL_1_xor54 = b_count_0_pad ^ state_1_pad;
  assign AXI4ToTL_1_xor26 = w_count_8_pad ^ AXI4ToTL_1_xor54;
  assign AXI4ToTL_1_xor12 = AXI4ToTL_1_xor25 ^ AXI4ToTL_1_xor26;
  assign AXI4ToTL_1_xor5 = AXI4ToTL_1_xor11 ^ AXI4ToTL_1_xor12;
  assign AXI4ToTL_1_xor27 = state_0_pad ^ w_count_15_pad;
  assign AXI4ToTL_1_xor28 = b_count_12_pad ^ w_count_11_pad;
  assign AXI4ToTL_1_xor13 = AXI4ToTL_1_xor27 ^ AXI4ToTL_1_xor28;
  assign AXI4ToTL_1_xor29 = b_count_9_pad ^ w_count_13_pad;
  assign AXI4ToTL_1_xor62 = b_count_15_pad ^ w_count_0_pad;
  assign AXI4ToTL_1_xor30 = w_count_5_pad ^ AXI4ToTL_1_xor62;
  assign AXI4ToTL_1_xor14 = AXI4ToTL_1_xor29 ^ AXI4ToTL_1_xor30;
  assign AXI4ToTL_1_xor6 = AXI4ToTL_1_xor13 ^ AXI4ToTL_1_xor14;
  assign AXI4ToTL_1_xor2 = AXI4ToTL_1_xor5 ^ AXI4ToTL_1_xor6;
  assign AXI4ToTL_1_xor0 = AXI4ToTL_1_xor1 ^ AXI4ToTL_1_xor2;
  assign deq_sum = AXI4ToTL_1_covSum + deq_io_covSum;
  assign q_b_deq_sum = deq_sum + q_b_deq_io_covSum;
  assign io_covSum = q_b_deq_sum;
  assign deq_metaReset = metaReset;
  assign q_b_deq_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_0 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[0]) begin
      r_count_0 <= _r_count_0_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_1 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[1]) begin
      r_count_1 <= _r_count_1_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_2 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[2]) begin
      r_count_2 <= _r_count_2_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_3 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[3]) begin
      r_count_3 <= _r_count_3_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_4 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[4]) begin
      r_count_4 <= _r_count_4_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_5 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[5]) begin
      r_count_5 <= _r_count_5_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_6 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[6]) begin
      r_count_6 <= _r_count_6_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_7 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[7]) begin
      r_count_7 <= _r_count_7_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_8 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[8]) begin
      r_count_8 <= _r_count_8_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_9 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[9]) begin
      r_count_9 <= _r_count_9_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_10 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[10]) begin
      r_count_10 <= _r_count_10_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_11 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[11]) begin
      r_count_11 <= _r_count_11_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_12 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[12]) begin
      r_count_12 <= _r_count_12_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_13 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[13]) begin
      r_count_13 <= _r_count_13_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_14 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[14]) begin
      r_count_14 <= _r_count_14_T_1;
    end
    if (reset) begin // @[ToTL.scala 91:28]
      r_count_15 <= 2'h0; // @[ToTL.scala 91:28]
    end else if (_T_26 & r_sel[15]) begin
      r_count_15 <= _r_count_15_T_1;
    end
    if (reset) begin // @[Arbiter.scala 87:30]
      beatsLeft <= 8'h0; // @[Arbiter.scala 87:30]
    end else if (latch) begin
      if (earlyWinner_1) begin
        beatsLeft <= auto_in_aw_bits_len;
      end else begin
        beatsLeft <= 8'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      readys_mask <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (latch & |readys_valid) begin
      readys_mask <= _readys_mask_T_3;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_0 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[0]) begin
      w_count_0 <= _w_count_0_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_1 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[1]) begin
      w_count_1 <= _w_count_1_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_2 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[2]) begin
      w_count_2 <= _w_count_2_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_3 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[3]) begin
      w_count_3 <= _w_count_3_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_4 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[4]) begin
      w_count_4 <= _w_count_4_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_5 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[5]) begin
      w_count_5 <= _w_count_5_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_6 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[6]) begin
      w_count_6 <= _w_count_6_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_7 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[7]) begin
      w_count_7 <= _w_count_7_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_8 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[8]) begin
      w_count_8 <= _w_count_8_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_9 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[9]) begin
      w_count_9 <= _w_count_9_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_10 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[10]) begin
      w_count_10 <= _w_count_10_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_11 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[11]) begin
      w_count_11 <= _w_count_11_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_12 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[12]) begin
      w_count_12 <= _w_count_12_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_13 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[13]) begin
      w_count_13 <= _w_count_13_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_14 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[14]) begin
      w_count_14 <= _w_count_14_T_1;
    end
    if (reset) begin // @[ToTL.scala 124:28]
      w_count_15 <= 2'h0; // @[ToTL.scala 124:28]
    end else if (_T_92 & w_sel[15]) begin
      w_count_15 <= _w_count_15_T_1;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      state_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (idle) begin
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Edges.scala 228:27]
      d_last_counter <= 9'h0; // @[Edges.scala 228:27]
    end else if (_d_last_T) begin
      if (d_last_first) begin
        if (d_hasData) begin
          d_last_counter <= d_last_beats1_decode;
        end else begin
          d_last_counter <= 9'h0;
        end
      end else begin
        d_last_counter <= d_last_counter1;
      end
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_0 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[0]) begin
      b_count_0 <= _b_count_0_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_1 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[1]) begin
      b_count_1 <= _b_count_1_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_2 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[2]) begin
      b_count_2 <= _b_count_2_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_3 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[3]) begin
      b_count_3 <= _b_count_3_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_4 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[4]) begin
      b_count_4 <= _b_count_4_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_5 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[5]) begin
      b_count_5 <= _b_count_5_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_6 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[6]) begin
      b_count_6 <= _b_count_6_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_7 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[7]) begin
      b_count_7 <= _b_count_7_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_8 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[8]) begin
      b_count_8 <= _b_count_8_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_9 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[9]) begin
      b_count_9 <= _b_count_9_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_10 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[10]) begin
      b_count_10 <= _b_count_10_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_11 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[11]) begin
      b_count_11 <= _b_count_11_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_12 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[12]) begin
      b_count_12 <= _b_count_12_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_13 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[13]) begin
      b_count_13 <= _b_count_13_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_14 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[14]) begin
      b_count_14 <= _b_count_14_T_1;
    end
    if (reset) begin // @[ToTL.scala 186:28]
      b_count_15 <= 2'h0; // @[ToTL.scala 186:28]
    end else if (_T_209 & b_sel[15]) begin
      b_count_15 <= _b_count_15_T_1;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_in_ar_valid | r_size1 == _T_4) & ~reset) begin
          $fatal; // @[ToTL.scala 98:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_in_ar_valid | r_size1 == _T_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:98 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n"
            ); // @[ToTL.scala 98:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_in_aw_valid | w_size1 == _T_62) & _T_8) begin
          $fatal; // @[ToTL.scala 131:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~auto_in_aw_valid | w_size1 == _T_62)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:131 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n"
            ); // @[ToTL.scala 131:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_58 | auto_in_aw_bits_len == 8'h0 | auto_in_aw_bits_size == 3'h3) & _T_8) begin
          $fatal; // @[ToTL.scala 132:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(_T_58 | auto_in_aw_bits_len == 8'h0 | auto_in_aw_bits_size == 3'h3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToTL.scala:132 assert (!in.aw.valid || in.aw.bits.len === UInt(0) || in.aw.bits.size === UInt(log2Ceil(beatBytes))) // because aligned\n"
            ); // @[ToTL.scala 132:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & _T_8) begin
          $fatal; // @[Arbiter.scala 22:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~earlyWinner_0 | ~earlyWinner_1) & _T_8) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~earlyWinner_0 | ~earlyWinner_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(auto_in_ar_valid | w_out_valid) | (earlyWinner_0 | earlyWinner_1)) & _T_8) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~(auto_in_ar_valid | w_out_valid) | (earlyWinner_0 | earlyWinner_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_135 | _T_134) & _T_8) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(_T_135 | _T_134)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    AXI4ToTL_1_covState <= AXI4ToTL_1_xor0;
    if (AXI4ToTL_1_covMap_write_en & AXI4ToTL_1_covMap_write_mask) begin
      AXI4ToTL_1_covMap[AXI4ToTL_1_covMap_write_addr] <= AXI4ToTL_1_covMap_write_data; // @[Coverage map for AXI4ToTL_1]
    end
    if (!(AXI4ToTL_1_covMap_read_data | metaReset)) begin
      AXI4ToTL_1_covSum <= AXI4ToTL_1_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    AXI4ToTL_1_covMap[initvar] = 0; //_54[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_count_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  r_count_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  r_count_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  r_count_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_count_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  r_count_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  r_count_6 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  r_count_7 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  r_count_8 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  r_count_9 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  r_count_10 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  r_count_11 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  r_count_12 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  r_count_13 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  r_count_14 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  r_count_15 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  beatsLeft = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  readys_mask = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  state_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  w_count_0 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  w_count_1 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  w_count_2 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  w_count_3 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  w_count_4 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  w_count_5 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  w_count_6 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  w_count_7 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  w_count_8 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  w_count_9 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  w_count_10 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  w_count_11 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  w_count_12 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  w_count_13 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  w_count_14 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  w_count_15 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  state_1 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  d_last_counter = _RAND_36[8:0];
  _RAND_37 = {1{`RANDOM}};
  b_count_0 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  b_count_1 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  b_count_2 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  b_count_3 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  b_count_4 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  b_count_5 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  b_count_6 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  b_count_7 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  b_count_8 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  b_count_9 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  b_count_10 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  b_count_11 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  b_count_12 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  b_count_13 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  b_count_14 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  b_count_15 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  AXI4ToTL_1_covState = 0; //_53[6:0];
  _RAND_55 = {1{`RANDOM}};
  AXI4ToTL_1_covSum = 0; //_55[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QueueCompatibility_36(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_real_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_real_last,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  ram_real_last [0:1]; // @[Decoupled.scala 259:95]
  wire  ram_real_last_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_real_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_real_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_real_last_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_real_last_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_real_last_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_real_last_MPORT_en; // @[Decoupled.scala 259:95]
  reg  enq_ptr_value; // @[Counter.scala 62:40]
  reg  deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] QueueCompatibility_36_covSum;
  assign ram_real_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_real_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_real_last_io_deq_bits_MPORT_data = ram_real_last[ram_real_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_real_last_MPORT_data = io_enq_bits_real_last;
  assign ram_real_last_MPORT_addr = enq_ptr_value;
  assign ram_real_last_MPORT_mask = 1'h1;
  assign ram_real_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_real_last = ram_real_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign QueueCompatibility_36_covSum = 30'h0;
  assign io_covSum = QueueCompatibility_36_covSum;
  always @(posedge clock) begin
    if (ram_real_last_MPORT_en & ram_real_last_MPORT_mask) begin
      ram_real_last[ram_real_last_MPORT_addr] <= ram_real_last_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      enq_ptr_value <= enq_ptr_value + 1'h1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 1'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      deq_ptr_value <= deq_ptr_value + 1'h1;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_real_last[initvar] = _RAND_0[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4UserYanker_2(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input         auto_in_aw_bits_echo_real_last,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_b_bits_echo_real_last,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input         auto_in_ar_bits_echo_real_last,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_echo_real_last,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last,
  output [29:0] io_covSum
);
  wire  QueueCompatibility_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_1_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_1_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_2_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_2_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_3_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_3_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_4_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_4_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_5_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_5_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_6_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_6_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_7_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_7_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_8_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_8_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_9_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_9_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_10_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_10_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_11_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_11_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_12_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_12_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_13_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_13_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_14_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_14_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_15_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_15_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_16_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_16_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_17_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_17_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_18_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_18_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_19_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_19_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_20_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_20_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_21_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_21_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_22_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_22_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_23_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_23_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_24_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_24_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_25_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_25_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_26_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_26_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_27_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_27_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_28_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_28_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_29_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_29_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_30_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_30_io_covSum; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_clock; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_reset; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_enq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_enq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_enq_bits_real_last; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_deq_ready; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_deq_valid; // @[UserYanker.scala 47:17]
  wire  QueueCompatibility_31_io_deq_bits_real_last; // @[UserYanker.scala 47:17]
  wire [29:0] QueueCompatibility_31_io_covSum; // @[UserYanker.scala 47:17]
  wire  _ar_ready_WIRE_0 = QueueCompatibility_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _ar_ready_WIRE_1 = QueueCompatibility_1_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_1 = 4'h1 == auto_in_ar_bits_id ? _ar_ready_WIRE_1 : _ar_ready_WIRE_0; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_2 = QueueCompatibility_2_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_2 = 4'h2 == auto_in_ar_bits_id ? _ar_ready_WIRE_2 : _GEN_1; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_3 = QueueCompatibility_3_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_3 = 4'h3 == auto_in_ar_bits_id ? _ar_ready_WIRE_3 : _GEN_2; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_4 = QueueCompatibility_4_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_4 = 4'h4 == auto_in_ar_bits_id ? _ar_ready_WIRE_4 : _GEN_3; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_5 = QueueCompatibility_5_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_5 = 4'h5 == auto_in_ar_bits_id ? _ar_ready_WIRE_5 : _GEN_4; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_6 = QueueCompatibility_6_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_6 = 4'h6 == auto_in_ar_bits_id ? _ar_ready_WIRE_6 : _GEN_5; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_7 = QueueCompatibility_7_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_7 = 4'h7 == auto_in_ar_bits_id ? _ar_ready_WIRE_7 : _GEN_6; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_8 = QueueCompatibility_8_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_8 = 4'h8 == auto_in_ar_bits_id ? _ar_ready_WIRE_8 : _GEN_7; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_9 = QueueCompatibility_9_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_9 = 4'h9 == auto_in_ar_bits_id ? _ar_ready_WIRE_9 : _GEN_8; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_10 = QueueCompatibility_10_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_10 = 4'ha == auto_in_ar_bits_id ? _ar_ready_WIRE_10 : _GEN_9; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_11 = QueueCompatibility_11_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_11 = 4'hb == auto_in_ar_bits_id ? _ar_ready_WIRE_11 : _GEN_10; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_12 = QueueCompatibility_12_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_12 = 4'hc == auto_in_ar_bits_id ? _ar_ready_WIRE_12 : _GEN_11; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_13 = QueueCompatibility_13_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_13 = 4'hd == auto_in_ar_bits_id ? _ar_ready_WIRE_13 : _GEN_12; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_14 = QueueCompatibility_14_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_14 = 4'he == auto_in_ar_bits_id ? _ar_ready_WIRE_14 : _GEN_13; // @[UserYanker.scala 56:{36,36}]
  wire  _ar_ready_WIRE_15 = QueueCompatibility_15_io_enq_ready; // @[UserYanker.scala 55:{25,25}]
  wire  _GEN_15 = 4'hf == auto_in_ar_bits_id ? _ar_ready_WIRE_15 : _GEN_14; // @[UserYanker.scala 56:{36,36}]
  wire  _r_valid_WIRE_0 = QueueCompatibility_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _r_valid_WIRE_1 = QueueCompatibility_1_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_17 = 4'h1 == auto_out_r_bits_id ? _r_valid_WIRE_1 : _r_valid_WIRE_0; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_2 = QueueCompatibility_2_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_18 = 4'h2 == auto_out_r_bits_id ? _r_valid_WIRE_2 : _GEN_17; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_3 = QueueCompatibility_3_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_19 = 4'h3 == auto_out_r_bits_id ? _r_valid_WIRE_3 : _GEN_18; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_4 = QueueCompatibility_4_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_20 = 4'h4 == auto_out_r_bits_id ? _r_valid_WIRE_4 : _GEN_19; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_5 = QueueCompatibility_5_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_21 = 4'h5 == auto_out_r_bits_id ? _r_valid_WIRE_5 : _GEN_20; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_6 = QueueCompatibility_6_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_22 = 4'h6 == auto_out_r_bits_id ? _r_valid_WIRE_6 : _GEN_21; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_7 = QueueCompatibility_7_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_23 = 4'h7 == auto_out_r_bits_id ? _r_valid_WIRE_7 : _GEN_22; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_8 = QueueCompatibility_8_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_24 = 4'h8 == auto_out_r_bits_id ? _r_valid_WIRE_8 : _GEN_23; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_9 = QueueCompatibility_9_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_25 = 4'h9 == auto_out_r_bits_id ? _r_valid_WIRE_9 : _GEN_24; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_10 = QueueCompatibility_10_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_26 = 4'ha == auto_out_r_bits_id ? _r_valid_WIRE_10 : _GEN_25; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_11 = QueueCompatibility_11_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_27 = 4'hb == auto_out_r_bits_id ? _r_valid_WIRE_11 : _GEN_26; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_12 = QueueCompatibility_12_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_28 = 4'hc == auto_out_r_bits_id ? _r_valid_WIRE_12 : _GEN_27; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_13 = QueueCompatibility_13_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_29 = 4'hd == auto_out_r_bits_id ? _r_valid_WIRE_13 : _GEN_28; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_14 = QueueCompatibility_14_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_30 = 4'he == auto_out_r_bits_id ? _r_valid_WIRE_14 : _GEN_29; // @[UserYanker.scala 63:{28,28}]
  wire  _r_valid_WIRE_15 = QueueCompatibility_15_io_deq_valid; // @[UserYanker.scala 61:{24,24}]
  wire  _GEN_31 = 4'hf == auto_out_r_bits_id ? _r_valid_WIRE_15 : _GEN_30; // @[UserYanker.scala 63:{28,28}]
  wire  _T_3 = ~reset; // @[UserYanker.scala 63:14]
  wire  _r_bits_WIRE_0_real_last = QueueCompatibility_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _r_bits_WIRE_1_real_last = QueueCompatibility_1_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_33 = 4'h1 == auto_out_r_bits_id ? _r_bits_WIRE_1_real_last : _r_bits_WIRE_0_real_last; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_2_real_last = QueueCompatibility_2_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_34 = 4'h2 == auto_out_r_bits_id ? _r_bits_WIRE_2_real_last : _GEN_33; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_3_real_last = QueueCompatibility_3_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_35 = 4'h3 == auto_out_r_bits_id ? _r_bits_WIRE_3_real_last : _GEN_34; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_4_real_last = QueueCompatibility_4_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_36 = 4'h4 == auto_out_r_bits_id ? _r_bits_WIRE_4_real_last : _GEN_35; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_5_real_last = QueueCompatibility_5_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_37 = 4'h5 == auto_out_r_bits_id ? _r_bits_WIRE_5_real_last : _GEN_36; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_6_real_last = QueueCompatibility_6_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_38 = 4'h6 == auto_out_r_bits_id ? _r_bits_WIRE_6_real_last : _GEN_37; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_7_real_last = QueueCompatibility_7_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_39 = 4'h7 == auto_out_r_bits_id ? _r_bits_WIRE_7_real_last : _GEN_38; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_8_real_last = QueueCompatibility_8_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_40 = 4'h8 == auto_out_r_bits_id ? _r_bits_WIRE_8_real_last : _GEN_39; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_9_real_last = QueueCompatibility_9_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_41 = 4'h9 == auto_out_r_bits_id ? _r_bits_WIRE_9_real_last : _GEN_40; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_10_real_last = QueueCompatibility_10_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_42 = 4'ha == auto_out_r_bits_id ? _r_bits_WIRE_10_real_last : _GEN_41; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_11_real_last = QueueCompatibility_11_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_43 = 4'hb == auto_out_r_bits_id ? _r_bits_WIRE_11_real_last : _GEN_42; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_12_real_last = QueueCompatibility_12_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_44 = 4'hc == auto_out_r_bits_id ? _r_bits_WIRE_12_real_last : _GEN_43; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_13_real_last = QueueCompatibility_13_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_45 = 4'hd == auto_out_r_bits_id ? _r_bits_WIRE_13_real_last : _GEN_44; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_14_real_last = QueueCompatibility_14_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire  _GEN_46 = 4'he == auto_out_r_bits_id ? _r_bits_WIRE_14_real_last : _GEN_45; // @[BundleMap.scala 247:{19,19}]
  wire  _r_bits_WIRE_15_real_last = QueueCompatibility_15_io_deq_bits_real_last; // @[UserYanker.scala 62:{23,23}]
  wire [15:0] _arsel_T = 16'h1 << auto_in_ar_bits_id; // @[OneHot.scala 64:12]
  wire  arsel_0 = _arsel_T[0]; // @[UserYanker.scala 67:55]
  wire  arsel_1 = _arsel_T[1]; // @[UserYanker.scala 67:55]
  wire  arsel_2 = _arsel_T[2]; // @[UserYanker.scala 67:55]
  wire  arsel_3 = _arsel_T[3]; // @[UserYanker.scala 67:55]
  wire  arsel_4 = _arsel_T[4]; // @[UserYanker.scala 67:55]
  wire  arsel_5 = _arsel_T[5]; // @[UserYanker.scala 67:55]
  wire  arsel_6 = _arsel_T[6]; // @[UserYanker.scala 67:55]
  wire  arsel_7 = _arsel_T[7]; // @[UserYanker.scala 67:55]
  wire  arsel_8 = _arsel_T[8]; // @[UserYanker.scala 67:55]
  wire  arsel_9 = _arsel_T[9]; // @[UserYanker.scala 67:55]
  wire  arsel_10 = _arsel_T[10]; // @[UserYanker.scala 67:55]
  wire  arsel_11 = _arsel_T[11]; // @[UserYanker.scala 67:55]
  wire  arsel_12 = _arsel_T[12]; // @[UserYanker.scala 67:55]
  wire  arsel_13 = _arsel_T[13]; // @[UserYanker.scala 67:55]
  wire  arsel_14 = _arsel_T[14]; // @[UserYanker.scala 67:55]
  wire  arsel_15 = _arsel_T[15]; // @[UserYanker.scala 67:55]
  wire [15:0] _rsel_T = 16'h1 << auto_out_r_bits_id; // @[OneHot.scala 64:12]
  wire  rsel_0 = _rsel_T[0]; // @[UserYanker.scala 68:55]
  wire  rsel_1 = _rsel_T[1]; // @[UserYanker.scala 68:55]
  wire  rsel_2 = _rsel_T[2]; // @[UserYanker.scala 68:55]
  wire  rsel_3 = _rsel_T[3]; // @[UserYanker.scala 68:55]
  wire  rsel_4 = _rsel_T[4]; // @[UserYanker.scala 68:55]
  wire  rsel_5 = _rsel_T[5]; // @[UserYanker.scala 68:55]
  wire  rsel_6 = _rsel_T[6]; // @[UserYanker.scala 68:55]
  wire  rsel_7 = _rsel_T[7]; // @[UserYanker.scala 68:55]
  wire  rsel_8 = _rsel_T[8]; // @[UserYanker.scala 68:55]
  wire  rsel_9 = _rsel_T[9]; // @[UserYanker.scala 68:55]
  wire  rsel_10 = _rsel_T[10]; // @[UserYanker.scala 68:55]
  wire  rsel_11 = _rsel_T[11]; // @[UserYanker.scala 68:55]
  wire  rsel_12 = _rsel_T[12]; // @[UserYanker.scala 68:55]
  wire  rsel_13 = _rsel_T[13]; // @[UserYanker.scala 68:55]
  wire  rsel_14 = _rsel_T[14]; // @[UserYanker.scala 68:55]
  wire  rsel_15 = _rsel_T[15]; // @[UserYanker.scala 68:55]
  wire  _aw_ready_WIRE_0 = QueueCompatibility_16_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _aw_ready_WIRE_1 = QueueCompatibility_17_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_49 = 4'h1 == auto_in_aw_bits_id ? _aw_ready_WIRE_1 : _aw_ready_WIRE_0; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_2 = QueueCompatibility_18_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_50 = 4'h2 == auto_in_aw_bits_id ? _aw_ready_WIRE_2 : _GEN_49; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_3 = QueueCompatibility_19_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_51 = 4'h3 == auto_in_aw_bits_id ? _aw_ready_WIRE_3 : _GEN_50; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_4 = QueueCompatibility_20_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_52 = 4'h4 == auto_in_aw_bits_id ? _aw_ready_WIRE_4 : _GEN_51; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_5 = QueueCompatibility_21_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_53 = 4'h5 == auto_in_aw_bits_id ? _aw_ready_WIRE_5 : _GEN_52; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_6 = QueueCompatibility_22_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_54 = 4'h6 == auto_in_aw_bits_id ? _aw_ready_WIRE_6 : _GEN_53; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_7 = QueueCompatibility_23_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_55 = 4'h7 == auto_in_aw_bits_id ? _aw_ready_WIRE_7 : _GEN_54; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_8 = QueueCompatibility_24_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_56 = 4'h8 == auto_in_aw_bits_id ? _aw_ready_WIRE_8 : _GEN_55; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_9 = QueueCompatibility_25_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_57 = 4'h9 == auto_in_aw_bits_id ? _aw_ready_WIRE_9 : _GEN_56; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_10 = QueueCompatibility_26_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_58 = 4'ha == auto_in_aw_bits_id ? _aw_ready_WIRE_10 : _GEN_57; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_11 = QueueCompatibility_27_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_59 = 4'hb == auto_in_aw_bits_id ? _aw_ready_WIRE_11 : _GEN_58; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_12 = QueueCompatibility_28_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_60 = 4'hc == auto_in_aw_bits_id ? _aw_ready_WIRE_12 : _GEN_59; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_13 = QueueCompatibility_29_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_61 = 4'hd == auto_in_aw_bits_id ? _aw_ready_WIRE_13 : _GEN_60; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_14 = QueueCompatibility_30_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_62 = 4'he == auto_in_aw_bits_id ? _aw_ready_WIRE_14 : _GEN_61; // @[UserYanker.scala 77:{36,36}]
  wire  _aw_ready_WIRE_15 = QueueCompatibility_31_io_enq_ready; // @[UserYanker.scala 76:{25,25}]
  wire  _GEN_63 = 4'hf == auto_in_aw_bits_id ? _aw_ready_WIRE_15 : _GEN_62; // @[UserYanker.scala 77:{36,36}]
  wire  _b_valid_WIRE_0 = QueueCompatibility_16_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _b_valid_WIRE_1 = QueueCompatibility_17_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_65 = 4'h1 == auto_out_b_bits_id ? _b_valid_WIRE_1 : _b_valid_WIRE_0; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_2 = QueueCompatibility_18_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_66 = 4'h2 == auto_out_b_bits_id ? _b_valid_WIRE_2 : _GEN_65; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_3 = QueueCompatibility_19_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_67 = 4'h3 == auto_out_b_bits_id ? _b_valid_WIRE_3 : _GEN_66; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_4 = QueueCompatibility_20_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_68 = 4'h4 == auto_out_b_bits_id ? _b_valid_WIRE_4 : _GEN_67; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_5 = QueueCompatibility_21_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_69 = 4'h5 == auto_out_b_bits_id ? _b_valid_WIRE_5 : _GEN_68; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_6 = QueueCompatibility_22_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_70 = 4'h6 == auto_out_b_bits_id ? _b_valid_WIRE_6 : _GEN_69; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_7 = QueueCompatibility_23_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_71 = 4'h7 == auto_out_b_bits_id ? _b_valid_WIRE_7 : _GEN_70; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_8 = QueueCompatibility_24_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_72 = 4'h8 == auto_out_b_bits_id ? _b_valid_WIRE_8 : _GEN_71; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_9 = QueueCompatibility_25_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_73 = 4'h9 == auto_out_b_bits_id ? _b_valid_WIRE_9 : _GEN_72; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_10 = QueueCompatibility_26_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_74 = 4'ha == auto_out_b_bits_id ? _b_valid_WIRE_10 : _GEN_73; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_11 = QueueCompatibility_27_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_75 = 4'hb == auto_out_b_bits_id ? _b_valid_WIRE_11 : _GEN_74; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_12 = QueueCompatibility_28_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_76 = 4'hc == auto_out_b_bits_id ? _b_valid_WIRE_12 : _GEN_75; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_13 = QueueCompatibility_29_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_77 = 4'hd == auto_out_b_bits_id ? _b_valid_WIRE_13 : _GEN_76; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_14 = QueueCompatibility_30_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_78 = 4'he == auto_out_b_bits_id ? _b_valid_WIRE_14 : _GEN_77; // @[UserYanker.scala 84:{28,28}]
  wire  _b_valid_WIRE_15 = QueueCompatibility_31_io_deq_valid; // @[UserYanker.scala 82:{24,24}]
  wire  _GEN_79 = 4'hf == auto_out_b_bits_id ? _b_valid_WIRE_15 : _GEN_78; // @[UserYanker.scala 84:{28,28}]
  wire  _b_bits_WIRE_0_real_last = QueueCompatibility_16_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _b_bits_WIRE_1_real_last = QueueCompatibility_17_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_81 = 4'h1 == auto_out_b_bits_id ? _b_bits_WIRE_1_real_last : _b_bits_WIRE_0_real_last; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_2_real_last = QueueCompatibility_18_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_82 = 4'h2 == auto_out_b_bits_id ? _b_bits_WIRE_2_real_last : _GEN_81; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_3_real_last = QueueCompatibility_19_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_83 = 4'h3 == auto_out_b_bits_id ? _b_bits_WIRE_3_real_last : _GEN_82; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_4_real_last = QueueCompatibility_20_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_84 = 4'h4 == auto_out_b_bits_id ? _b_bits_WIRE_4_real_last : _GEN_83; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_5_real_last = QueueCompatibility_21_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_85 = 4'h5 == auto_out_b_bits_id ? _b_bits_WIRE_5_real_last : _GEN_84; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_6_real_last = QueueCompatibility_22_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_86 = 4'h6 == auto_out_b_bits_id ? _b_bits_WIRE_6_real_last : _GEN_85; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_7_real_last = QueueCompatibility_23_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_87 = 4'h7 == auto_out_b_bits_id ? _b_bits_WIRE_7_real_last : _GEN_86; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_8_real_last = QueueCompatibility_24_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_88 = 4'h8 == auto_out_b_bits_id ? _b_bits_WIRE_8_real_last : _GEN_87; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_9_real_last = QueueCompatibility_25_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_89 = 4'h9 == auto_out_b_bits_id ? _b_bits_WIRE_9_real_last : _GEN_88; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_10_real_last = QueueCompatibility_26_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_90 = 4'ha == auto_out_b_bits_id ? _b_bits_WIRE_10_real_last : _GEN_89; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_11_real_last = QueueCompatibility_27_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_91 = 4'hb == auto_out_b_bits_id ? _b_bits_WIRE_11_real_last : _GEN_90; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_12_real_last = QueueCompatibility_28_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_92 = 4'hc == auto_out_b_bits_id ? _b_bits_WIRE_12_real_last : _GEN_91; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_13_real_last = QueueCompatibility_29_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_93 = 4'hd == auto_out_b_bits_id ? _b_bits_WIRE_13_real_last : _GEN_92; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_14_real_last = QueueCompatibility_30_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire  _GEN_94 = 4'he == auto_out_b_bits_id ? _b_bits_WIRE_14_real_last : _GEN_93; // @[BundleMap.scala 247:{19,19}]
  wire  _b_bits_WIRE_15_real_last = QueueCompatibility_31_io_deq_bits_real_last; // @[UserYanker.scala 83:{23,23}]
  wire [15:0] _awsel_T = 16'h1 << auto_in_aw_bits_id; // @[OneHot.scala 64:12]
  wire  awsel_0 = _awsel_T[0]; // @[UserYanker.scala 88:55]
  wire  awsel_1 = _awsel_T[1]; // @[UserYanker.scala 88:55]
  wire  awsel_2 = _awsel_T[2]; // @[UserYanker.scala 88:55]
  wire  awsel_3 = _awsel_T[3]; // @[UserYanker.scala 88:55]
  wire  awsel_4 = _awsel_T[4]; // @[UserYanker.scala 88:55]
  wire  awsel_5 = _awsel_T[5]; // @[UserYanker.scala 88:55]
  wire  awsel_6 = _awsel_T[6]; // @[UserYanker.scala 88:55]
  wire  awsel_7 = _awsel_T[7]; // @[UserYanker.scala 88:55]
  wire  awsel_8 = _awsel_T[8]; // @[UserYanker.scala 88:55]
  wire  awsel_9 = _awsel_T[9]; // @[UserYanker.scala 88:55]
  wire  awsel_10 = _awsel_T[10]; // @[UserYanker.scala 88:55]
  wire  awsel_11 = _awsel_T[11]; // @[UserYanker.scala 88:55]
  wire  awsel_12 = _awsel_T[12]; // @[UserYanker.scala 88:55]
  wire  awsel_13 = _awsel_T[13]; // @[UserYanker.scala 88:55]
  wire  awsel_14 = _awsel_T[14]; // @[UserYanker.scala 88:55]
  wire  awsel_15 = _awsel_T[15]; // @[UserYanker.scala 88:55]
  wire [15:0] _bsel_T = 16'h1 << auto_out_b_bits_id; // @[OneHot.scala 64:12]
  wire  bsel_0 = _bsel_T[0]; // @[UserYanker.scala 89:55]
  wire  bsel_1 = _bsel_T[1]; // @[UserYanker.scala 89:55]
  wire  bsel_2 = _bsel_T[2]; // @[UserYanker.scala 89:55]
  wire  bsel_3 = _bsel_T[3]; // @[UserYanker.scala 89:55]
  wire  bsel_4 = _bsel_T[4]; // @[UserYanker.scala 89:55]
  wire  bsel_5 = _bsel_T[5]; // @[UserYanker.scala 89:55]
  wire  bsel_6 = _bsel_T[6]; // @[UserYanker.scala 89:55]
  wire  bsel_7 = _bsel_T[7]; // @[UserYanker.scala 89:55]
  wire  bsel_8 = _bsel_T[8]; // @[UserYanker.scala 89:55]
  wire  bsel_9 = _bsel_T[9]; // @[UserYanker.scala 89:55]
  wire  bsel_10 = _bsel_T[10]; // @[UserYanker.scala 89:55]
  wire  bsel_11 = _bsel_T[11]; // @[UserYanker.scala 89:55]
  wire  bsel_12 = _bsel_T[12]; // @[UserYanker.scala 89:55]
  wire  bsel_13 = _bsel_T[13]; // @[UserYanker.scala 89:55]
  wire  bsel_14 = _bsel_T[14]; // @[UserYanker.scala 89:55]
  wire  bsel_15 = _bsel_T[15]; // @[UserYanker.scala 89:55]
  wire [29:0] AXI4UserYanker_2_covSum;
  wire [29:0] QueueCompatibility_19_sum;
  wire [29:0] QueueCompatibility_14_sum;
  wire [29:0] QueueCompatibility_12_sum;
  wire [29:0] QueueCompatibility_9_sum;
  wire [29:0] QueueCompatibility_31_sum;
  wire [29:0] QueueCompatibility_29_sum;
  wire [29:0] QueueCompatibility_3_sum;
  wire [29:0] QueueCompatibility_26_sum;
  wire [29:0] QueueCompatibility_28_sum;
  wire [29:0] QueueCompatibility_16_sum;
  wire [29:0] QueueCompatibility_8_sum;
  wire [29:0] QueueCompatibility_sum;
  wire [29:0] QueueCompatibility_5_sum;
  wire [29:0] QueueCompatibility_17_sum;
  wire [29:0] QueueCompatibility_27_sum;
  wire [29:0] QueueCompatibility_24_sum;
  wire [29:0] QueueCompatibility_6_sum;
  wire [29:0] QueueCompatibility_22_sum;
  wire [29:0] QueueCompatibility_18_sum;
  wire [29:0] QueueCompatibility_13_sum;
  wire [29:0] QueueCompatibility_11_sum;
  wire [29:0] QueueCompatibility_1_sum;
  wire [29:0] QueueCompatibility_21_sum;
  wire [29:0] QueueCompatibility_30_sum;
  wire [29:0] QueueCompatibility_25_sum;
  wire [29:0] QueueCompatibility_7_sum;
  wire [29:0] QueueCompatibility_20_sum;
  wire [29:0] QueueCompatibility_4_sum;
  wire [29:0] QueueCompatibility_10_sum;
  wire [29:0] QueueCompatibility_23_sum;
  wire [29:0] QueueCompatibility_2_sum;
  wire [29:0] QueueCompatibility_15_sum;
  QueueCompatibility_36 QueueCompatibility ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_clock),
    .reset(QueueCompatibility_reset),
    .io_enq_ready(QueueCompatibility_io_enq_ready),
    .io_enq_valid(QueueCompatibility_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_io_deq_ready),
    .io_deq_valid(QueueCompatibility_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_1 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_1_clock),
    .reset(QueueCompatibility_1_reset),
    .io_enq_ready(QueueCompatibility_1_io_enq_ready),
    .io_enq_valid(QueueCompatibility_1_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_1_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_1_io_deq_ready),
    .io_deq_valid(QueueCompatibility_1_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_1_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_1_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_2 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_2_clock),
    .reset(QueueCompatibility_2_reset),
    .io_enq_ready(QueueCompatibility_2_io_enq_ready),
    .io_enq_valid(QueueCompatibility_2_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_2_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_2_io_deq_ready),
    .io_deq_valid(QueueCompatibility_2_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_2_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_2_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_3 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_3_clock),
    .reset(QueueCompatibility_3_reset),
    .io_enq_ready(QueueCompatibility_3_io_enq_ready),
    .io_enq_valid(QueueCompatibility_3_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_3_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_3_io_deq_ready),
    .io_deq_valid(QueueCompatibility_3_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_3_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_3_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_4 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_4_clock),
    .reset(QueueCompatibility_4_reset),
    .io_enq_ready(QueueCompatibility_4_io_enq_ready),
    .io_enq_valid(QueueCompatibility_4_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_4_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_4_io_deq_ready),
    .io_deq_valid(QueueCompatibility_4_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_4_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_4_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_5 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_5_clock),
    .reset(QueueCompatibility_5_reset),
    .io_enq_ready(QueueCompatibility_5_io_enq_ready),
    .io_enq_valid(QueueCompatibility_5_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_5_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_5_io_deq_ready),
    .io_deq_valid(QueueCompatibility_5_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_5_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_5_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_6 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_6_clock),
    .reset(QueueCompatibility_6_reset),
    .io_enq_ready(QueueCompatibility_6_io_enq_ready),
    .io_enq_valid(QueueCompatibility_6_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_6_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_6_io_deq_ready),
    .io_deq_valid(QueueCompatibility_6_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_6_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_6_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_7 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_7_clock),
    .reset(QueueCompatibility_7_reset),
    .io_enq_ready(QueueCompatibility_7_io_enq_ready),
    .io_enq_valid(QueueCompatibility_7_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_7_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_7_io_deq_ready),
    .io_deq_valid(QueueCompatibility_7_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_7_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_7_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_8 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_8_clock),
    .reset(QueueCompatibility_8_reset),
    .io_enq_ready(QueueCompatibility_8_io_enq_ready),
    .io_enq_valid(QueueCompatibility_8_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_8_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_8_io_deq_ready),
    .io_deq_valid(QueueCompatibility_8_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_8_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_8_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_9 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_9_clock),
    .reset(QueueCompatibility_9_reset),
    .io_enq_ready(QueueCompatibility_9_io_enq_ready),
    .io_enq_valid(QueueCompatibility_9_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_9_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_9_io_deq_ready),
    .io_deq_valid(QueueCompatibility_9_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_9_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_9_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_10 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_10_clock),
    .reset(QueueCompatibility_10_reset),
    .io_enq_ready(QueueCompatibility_10_io_enq_ready),
    .io_enq_valid(QueueCompatibility_10_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_10_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_10_io_deq_ready),
    .io_deq_valid(QueueCompatibility_10_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_10_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_10_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_11 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_11_clock),
    .reset(QueueCompatibility_11_reset),
    .io_enq_ready(QueueCompatibility_11_io_enq_ready),
    .io_enq_valid(QueueCompatibility_11_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_11_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_11_io_deq_ready),
    .io_deq_valid(QueueCompatibility_11_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_11_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_11_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_12 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_12_clock),
    .reset(QueueCompatibility_12_reset),
    .io_enq_ready(QueueCompatibility_12_io_enq_ready),
    .io_enq_valid(QueueCompatibility_12_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_12_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_12_io_deq_ready),
    .io_deq_valid(QueueCompatibility_12_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_12_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_12_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_13 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_13_clock),
    .reset(QueueCompatibility_13_reset),
    .io_enq_ready(QueueCompatibility_13_io_enq_ready),
    .io_enq_valid(QueueCompatibility_13_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_13_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_13_io_deq_ready),
    .io_deq_valid(QueueCompatibility_13_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_13_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_13_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_14 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_14_clock),
    .reset(QueueCompatibility_14_reset),
    .io_enq_ready(QueueCompatibility_14_io_enq_ready),
    .io_enq_valid(QueueCompatibility_14_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_14_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_14_io_deq_ready),
    .io_deq_valid(QueueCompatibility_14_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_14_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_14_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_15 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_15_clock),
    .reset(QueueCompatibility_15_reset),
    .io_enq_ready(QueueCompatibility_15_io_enq_ready),
    .io_enq_valid(QueueCompatibility_15_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_15_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_15_io_deq_ready),
    .io_deq_valid(QueueCompatibility_15_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_15_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_15_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_16 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_16_clock),
    .reset(QueueCompatibility_16_reset),
    .io_enq_ready(QueueCompatibility_16_io_enq_ready),
    .io_enq_valid(QueueCompatibility_16_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_16_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_16_io_deq_ready),
    .io_deq_valid(QueueCompatibility_16_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_16_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_16_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_17 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_17_clock),
    .reset(QueueCompatibility_17_reset),
    .io_enq_ready(QueueCompatibility_17_io_enq_ready),
    .io_enq_valid(QueueCompatibility_17_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_17_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_17_io_deq_ready),
    .io_deq_valid(QueueCompatibility_17_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_17_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_17_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_18 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_18_clock),
    .reset(QueueCompatibility_18_reset),
    .io_enq_ready(QueueCompatibility_18_io_enq_ready),
    .io_enq_valid(QueueCompatibility_18_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_18_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_18_io_deq_ready),
    .io_deq_valid(QueueCompatibility_18_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_18_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_18_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_19 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_19_clock),
    .reset(QueueCompatibility_19_reset),
    .io_enq_ready(QueueCompatibility_19_io_enq_ready),
    .io_enq_valid(QueueCompatibility_19_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_19_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_19_io_deq_ready),
    .io_deq_valid(QueueCompatibility_19_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_19_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_19_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_20 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_20_clock),
    .reset(QueueCompatibility_20_reset),
    .io_enq_ready(QueueCompatibility_20_io_enq_ready),
    .io_enq_valid(QueueCompatibility_20_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_20_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_20_io_deq_ready),
    .io_deq_valid(QueueCompatibility_20_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_20_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_20_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_21 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_21_clock),
    .reset(QueueCompatibility_21_reset),
    .io_enq_ready(QueueCompatibility_21_io_enq_ready),
    .io_enq_valid(QueueCompatibility_21_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_21_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_21_io_deq_ready),
    .io_deq_valid(QueueCompatibility_21_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_21_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_21_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_22 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_22_clock),
    .reset(QueueCompatibility_22_reset),
    .io_enq_ready(QueueCompatibility_22_io_enq_ready),
    .io_enq_valid(QueueCompatibility_22_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_22_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_22_io_deq_ready),
    .io_deq_valid(QueueCompatibility_22_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_22_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_22_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_23 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_23_clock),
    .reset(QueueCompatibility_23_reset),
    .io_enq_ready(QueueCompatibility_23_io_enq_ready),
    .io_enq_valid(QueueCompatibility_23_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_23_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_23_io_deq_ready),
    .io_deq_valid(QueueCompatibility_23_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_23_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_23_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_24 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_24_clock),
    .reset(QueueCompatibility_24_reset),
    .io_enq_ready(QueueCompatibility_24_io_enq_ready),
    .io_enq_valid(QueueCompatibility_24_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_24_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_24_io_deq_ready),
    .io_deq_valid(QueueCompatibility_24_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_24_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_24_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_25 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_25_clock),
    .reset(QueueCompatibility_25_reset),
    .io_enq_ready(QueueCompatibility_25_io_enq_ready),
    .io_enq_valid(QueueCompatibility_25_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_25_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_25_io_deq_ready),
    .io_deq_valid(QueueCompatibility_25_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_25_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_25_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_26 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_26_clock),
    .reset(QueueCompatibility_26_reset),
    .io_enq_ready(QueueCompatibility_26_io_enq_ready),
    .io_enq_valid(QueueCompatibility_26_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_26_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_26_io_deq_ready),
    .io_deq_valid(QueueCompatibility_26_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_26_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_26_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_27 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_27_clock),
    .reset(QueueCompatibility_27_reset),
    .io_enq_ready(QueueCompatibility_27_io_enq_ready),
    .io_enq_valid(QueueCompatibility_27_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_27_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_27_io_deq_ready),
    .io_deq_valid(QueueCompatibility_27_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_27_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_27_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_28 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_28_clock),
    .reset(QueueCompatibility_28_reset),
    .io_enq_ready(QueueCompatibility_28_io_enq_ready),
    .io_enq_valid(QueueCompatibility_28_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_28_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_28_io_deq_ready),
    .io_deq_valid(QueueCompatibility_28_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_28_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_28_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_29 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_29_clock),
    .reset(QueueCompatibility_29_reset),
    .io_enq_ready(QueueCompatibility_29_io_enq_ready),
    .io_enq_valid(QueueCompatibility_29_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_29_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_29_io_deq_ready),
    .io_deq_valid(QueueCompatibility_29_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_29_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_29_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_30 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_30_clock),
    .reset(QueueCompatibility_30_reset),
    .io_enq_ready(QueueCompatibility_30_io_enq_ready),
    .io_enq_valid(QueueCompatibility_30_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_30_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_30_io_deq_ready),
    .io_deq_valid(QueueCompatibility_30_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_30_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_30_io_covSum)
  );
  QueueCompatibility_36 QueueCompatibility_31 ( // @[UserYanker.scala 47:17]
    .clock(QueueCompatibility_31_clock),
    .reset(QueueCompatibility_31_reset),
    .io_enq_ready(QueueCompatibility_31_io_enq_ready),
    .io_enq_valid(QueueCompatibility_31_io_enq_valid),
    .io_enq_bits_real_last(QueueCompatibility_31_io_enq_bits_real_last),
    .io_deq_ready(QueueCompatibility_31_io_deq_ready),
    .io_deq_valid(QueueCompatibility_31_io_deq_valid),
    .io_deq_bits_real_last(QueueCompatibility_31_io_deq_bits_real_last),
    .io_covSum(QueueCompatibility_31_io_covSum)
  );
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_63; // @[UserYanker.scala 77:36]
  assign auto_in_w_ready = auto_out_w_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_echo_real_last = 4'hf == auto_out_b_bits_id ? _b_bits_WIRE_15_real_last : _GEN_94; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_15; // @[UserYanker.scala 56:36]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_echo_real_last = 4'hf == auto_out_r_bits_id ? _r_bits_WIRE_15_real_last : _GEN_46; // @[BundleMap.scala 247:{19,19}]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_63; // @[UserYanker.scala 78:36]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_valid = auto_in_w_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_15; // @[UserYanker.scala 57:36]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_clock = clock;
  assign QueueCompatibility_reset = reset;
  assign QueueCompatibility_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_0; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_0 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_1_clock = clock;
  assign QueueCompatibility_1_reset = reset;
  assign QueueCompatibility_1_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_1; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_1_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_1_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_1 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_2_clock = clock;
  assign QueueCompatibility_2_reset = reset;
  assign QueueCompatibility_2_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_2; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_2_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_2_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_2 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_3_clock = clock;
  assign QueueCompatibility_3_reset = reset;
  assign QueueCompatibility_3_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_3; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_3_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_3_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_3 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_4_clock = clock;
  assign QueueCompatibility_4_reset = reset;
  assign QueueCompatibility_4_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_4; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_4_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_4_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_4 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_5_clock = clock;
  assign QueueCompatibility_5_reset = reset;
  assign QueueCompatibility_5_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_5; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_5_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_5_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_5 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_6_clock = clock;
  assign QueueCompatibility_6_reset = reset;
  assign QueueCompatibility_6_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_6; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_6_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_6_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_6 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_7_clock = clock;
  assign QueueCompatibility_7_reset = reset;
  assign QueueCompatibility_7_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_7; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_7_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_7_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_7 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_8_clock = clock;
  assign QueueCompatibility_8_reset = reset;
  assign QueueCompatibility_8_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_8; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_8_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_8_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_8 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_9_clock = clock;
  assign QueueCompatibility_9_reset = reset;
  assign QueueCompatibility_9_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_9; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_9_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_9_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_9 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_10_clock = clock;
  assign QueueCompatibility_10_reset = reset;
  assign QueueCompatibility_10_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_10; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_10_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_10_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_10 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_11_clock = clock;
  assign QueueCompatibility_11_reset = reset;
  assign QueueCompatibility_11_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_11; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_11_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_11_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_11 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_12_clock = clock;
  assign QueueCompatibility_12_reset = reset;
  assign QueueCompatibility_12_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_12; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_12_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_12_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_12 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_13_clock = clock;
  assign QueueCompatibility_13_reset = reset;
  assign QueueCompatibility_13_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_13; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_13_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_13_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_13 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_14_clock = clock;
  assign QueueCompatibility_14_reset = reset;
  assign QueueCompatibility_14_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_14; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_14_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_14_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_14 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_15_clock = clock;
  assign QueueCompatibility_15_reset = reset;
  assign QueueCompatibility_15_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_15; // @[UserYanker.scala 71:53]
  assign QueueCompatibility_15_io_enq_bits_real_last = auto_in_ar_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_15_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_15 & auto_out_r_bits_last; // @[UserYanker.scala 70:58]
  assign QueueCompatibility_16_clock = clock;
  assign QueueCompatibility_16_reset = reset;
  assign QueueCompatibility_16_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_0; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_16_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_16_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_0; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_17_clock = clock;
  assign QueueCompatibility_17_reset = reset;
  assign QueueCompatibility_17_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_1; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_17_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_17_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_1; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_18_clock = clock;
  assign QueueCompatibility_18_reset = reset;
  assign QueueCompatibility_18_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_2; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_18_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_18_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_2; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_19_clock = clock;
  assign QueueCompatibility_19_reset = reset;
  assign QueueCompatibility_19_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_3; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_19_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_19_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_3; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_20_clock = clock;
  assign QueueCompatibility_20_reset = reset;
  assign QueueCompatibility_20_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_4; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_20_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_20_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_4; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_21_clock = clock;
  assign QueueCompatibility_21_reset = reset;
  assign QueueCompatibility_21_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_5; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_21_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_21_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_5; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_22_clock = clock;
  assign QueueCompatibility_22_reset = reset;
  assign QueueCompatibility_22_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_6; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_22_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_22_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_6; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_23_clock = clock;
  assign QueueCompatibility_23_reset = reset;
  assign QueueCompatibility_23_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_7; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_23_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_23_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_7; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_24_clock = clock;
  assign QueueCompatibility_24_reset = reset;
  assign QueueCompatibility_24_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_8; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_24_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_24_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_8; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_25_clock = clock;
  assign QueueCompatibility_25_reset = reset;
  assign QueueCompatibility_25_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_9; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_25_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_25_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_9; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_26_clock = clock;
  assign QueueCompatibility_26_reset = reset;
  assign QueueCompatibility_26_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_10; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_26_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_26_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_10; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_27_clock = clock;
  assign QueueCompatibility_27_reset = reset;
  assign QueueCompatibility_27_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_11; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_27_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_27_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_11; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_28_clock = clock;
  assign QueueCompatibility_28_reset = reset;
  assign QueueCompatibility_28_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_12; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_28_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_28_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_12; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_29_clock = clock;
  assign QueueCompatibility_29_reset = reset;
  assign QueueCompatibility_29_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_13; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_29_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_29_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_13; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_30_clock = clock;
  assign QueueCompatibility_30_reset = reset;
  assign QueueCompatibility_30_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_14; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_30_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_30_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_14; // @[UserYanker.scala 91:53]
  assign QueueCompatibility_31_clock = clock;
  assign QueueCompatibility_31_reset = reset;
  assign QueueCompatibility_31_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_15; // @[UserYanker.scala 92:53]
  assign QueueCompatibility_31_io_enq_bits_real_last = auto_in_aw_bits_echo_real_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign QueueCompatibility_31_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_15; // @[UserYanker.scala 91:53]
  assign AXI4UserYanker_2_covSum = 30'h0;
  assign QueueCompatibility_19_sum = AXI4UserYanker_2_covSum + QueueCompatibility_19_io_covSum;
  assign QueueCompatibility_14_sum = QueueCompatibility_19_sum + QueueCompatibility_14_io_covSum;
  assign QueueCompatibility_12_sum = QueueCompatibility_14_sum + QueueCompatibility_12_io_covSum;
  assign QueueCompatibility_9_sum = QueueCompatibility_12_sum + QueueCompatibility_9_io_covSum;
  assign QueueCompatibility_31_sum = QueueCompatibility_9_sum + QueueCompatibility_31_io_covSum;
  assign QueueCompatibility_29_sum = QueueCompatibility_31_sum + QueueCompatibility_29_io_covSum;
  assign QueueCompatibility_3_sum = QueueCompatibility_29_sum + QueueCompatibility_3_io_covSum;
  assign QueueCompatibility_26_sum = QueueCompatibility_3_sum + QueueCompatibility_26_io_covSum;
  assign QueueCompatibility_28_sum = QueueCompatibility_26_sum + QueueCompatibility_28_io_covSum;
  assign QueueCompatibility_16_sum = QueueCompatibility_28_sum + QueueCompatibility_16_io_covSum;
  assign QueueCompatibility_8_sum = QueueCompatibility_16_sum + QueueCompatibility_8_io_covSum;
  assign QueueCompatibility_sum = QueueCompatibility_8_sum + QueueCompatibility_io_covSum;
  assign QueueCompatibility_5_sum = QueueCompatibility_sum + QueueCompatibility_5_io_covSum;
  assign QueueCompatibility_17_sum = QueueCompatibility_5_sum + QueueCompatibility_17_io_covSum;
  assign QueueCompatibility_27_sum = QueueCompatibility_17_sum + QueueCompatibility_27_io_covSum;
  assign QueueCompatibility_24_sum = QueueCompatibility_27_sum + QueueCompatibility_24_io_covSum;
  assign QueueCompatibility_6_sum = QueueCompatibility_24_sum + QueueCompatibility_6_io_covSum;
  assign QueueCompatibility_22_sum = QueueCompatibility_6_sum + QueueCompatibility_22_io_covSum;
  assign QueueCompatibility_18_sum = QueueCompatibility_22_sum + QueueCompatibility_18_io_covSum;
  assign QueueCompatibility_13_sum = QueueCompatibility_18_sum + QueueCompatibility_13_io_covSum;
  assign QueueCompatibility_11_sum = QueueCompatibility_13_sum + QueueCompatibility_11_io_covSum;
  assign QueueCompatibility_1_sum = QueueCompatibility_11_sum + QueueCompatibility_1_io_covSum;
  assign QueueCompatibility_21_sum = QueueCompatibility_1_sum + QueueCompatibility_21_io_covSum;
  assign QueueCompatibility_30_sum = QueueCompatibility_21_sum + QueueCompatibility_30_io_covSum;
  assign QueueCompatibility_25_sum = QueueCompatibility_30_sum + QueueCompatibility_25_io_covSum;
  assign QueueCompatibility_7_sum = QueueCompatibility_25_sum + QueueCompatibility_7_io_covSum;
  assign QueueCompatibility_20_sum = QueueCompatibility_7_sum + QueueCompatibility_20_io_covSum;
  assign QueueCompatibility_4_sum = QueueCompatibility_20_sum + QueueCompatibility_4_io_covSum;
  assign QueueCompatibility_10_sum = QueueCompatibility_4_sum + QueueCompatibility_10_io_covSum;
  assign QueueCompatibility_23_sum = QueueCompatibility_10_sum + QueueCompatibility_23_io_covSum;
  assign QueueCompatibility_2_sum = QueueCompatibility_23_sum + QueueCompatibility_2_io_covSum;
  assign QueueCompatibility_15_sum = QueueCompatibility_2_sum + QueueCompatibility_15_io_covSum;
  assign io_covSum = QueueCompatibility_15_sum;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_r_valid | _GEN_31) & ~reset) begin
          $fatal; // @[UserYanker.scala 63:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_out_r_valid | _GEN_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:63 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 63:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~auto_out_b_valid | _GEN_79) & _T_3) begin
          $fatal; // @[UserYanker.scala 84:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~auto_out_b_valid | _GEN_79)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:84 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"
            ); // @[UserYanker.scala 84:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_28(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input  [3:0]  io_enq_bits_cache,
  input  [2:0]  io_enq_bits_prot,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output [3:0]  io_deq_bits_cache,
  output [2:0]  io_deq_bits_prot,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_id_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 259:95]
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_len [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_len_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_burst [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_burst_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_burst_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_cache [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_cache_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_cache_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_cache_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_cache_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] ram_prot [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_prot_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_prot_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [2:0] ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_prot_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_prot_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_17 = io_deq_ready ? 1'h0 : _do_enq_T; // @[Decoupled.scala 304:{26,35}]
  wire  do_enq = empty ? _GEN_17 : _do_enq_T; // @[Decoupled.scala 301:17]
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[Decoupled.scala 301:17 303:14]
  reg  Queue_28_covState; // @[Register tracking Queue_28 state]
  reg  Queue_28_covMap [0:1]; // @[Coverage map for Queue_28]
  wire  Queue_28_covMap_read_en; // @[Coverage map for Queue_28]
  wire  Queue_28_covMap_read_addr; // @[Coverage map for Queue_28]
  wire  Queue_28_covMap_read_data; // @[Coverage map for Queue_28]
  wire  Queue_28_covMap_write_data; // @[Coverage map for Queue_28]
  wire  Queue_28_covMap_write_addr; // @[Coverage map for Queue_28]
  wire  Queue_28_covMap_write_mask; // @[Coverage map for Queue_28]
  wire  Queue_28_covMap_write_en; // @[Coverage map for Queue_28]
  reg [29:0] Queue_28_covSum; // @[Sum of coverage map]
  wire  maybe_full_shl;
  wire  maybe_full_pad;
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_cache_io_deq_bits_MPORT_en = 1'h1;
  assign ram_cache_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_cache_io_deq_bits_MPORT_data = ram_cache[ram_cache_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_cache_MPORT_data = io_enq_bits_cache;
  assign ram_cache_MPORT_addr = 1'h0;
  assign ram_cache_MPORT_mask = 1'h1;
  assign ram_cache_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_prot_io_deq_bits_MPORT_en = 1'h1;
  assign ram_prot_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_prot_io_deq_bits_MPORT_data = ram_prot[ram_prot_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_prot_MPORT_data = io_enq_bits_prot;
  assign ram_prot_MPORT_addr = 1'h0;
  assign ram_prot_MPORT_mask = 1'h1;
  assign ram_prot_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[Decoupled.scala 288:16 300:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_burst = empty ? io_enq_bits_burst : ram_burst_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_cache = empty ? io_enq_bits_cache : ram_cache_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign io_deq_bits_prot = empty ? io_enq_bits_prot : ram_prot_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17 301:17 302:19]
  assign Queue_28_covMap_read_en = 1'h1;
  assign Queue_28_covMap_read_addr = Queue_28_covState;
  assign Queue_28_covMap_read_data = Queue_28_covMap[Queue_28_covMap_read_addr]; // @[Coverage map for Queue_28]
  assign Queue_28_covMap_write_data = 1'h1;
  assign Queue_28_covMap_write_addr = Queue_28_covState;
  assign Queue_28_covMap_write_mask = 1'h1;
  assign Queue_28_covMap_write_en = ~metaReset;
  assign maybe_full_shl = maybe_full;
  assign maybe_full_pad = maybe_full_shl;
  assign io_covSum = Queue_28_covSum;
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_cache_MPORT_en & ram_cache_MPORT_mask) begin
      ram_cache[ram_cache_MPORT_addr] <= ram_cache_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_prot_MPORT_en & ram_prot_MPORT_mask) begin
      ram_prot[ram_prot_MPORT_addr] <= ram_prot_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      if (empty) begin
        if (io_deq_ready) begin
          maybe_full <= 1'h0;
        end else begin
          maybe_full <= _do_enq_T;
        end
      end else begin
        maybe_full <= _do_enq_T;
      end
    end
    Queue_28_covState <= maybe_full_pad;
    if (Queue_28_covMap_write_en & Queue_28_covMap_write_mask) begin
      Queue_28_covMap[Queue_28_covMap_write_addr] <= Queue_28_covMap_write_data; // @[Coverage map for Queue_28]
    end
    if (!(Queue_28_covMap_read_data | metaReset)) begin
      Queue_28_covSum <= Queue_28_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = _RAND_6[2:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    Queue_28_covMap[initvar] = 0; //_9[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  Queue_28_covState = 0; //_8[0:0];
  _RAND_10 = {1{`RANDOM}};
  Queue_28_covSum = 0; //_10[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4Fragmenter_1(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output        auto_out_aw_bits_echo_real_last,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_b_bits_echo_real_last,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output        auto_out_ar_bits_echo_real_last,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_echo_real_last,
  input         auto_out_r_bits_last,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_25;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  wire  deq_clock; // @[Decoupled.scala 361:21]
  wire  deq_reset; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] deq_io_enq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] deq_io_enq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] deq_io_enq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] deq_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] deq_io_enq_bits_burst; // @[Decoupled.scala 361:21]
  wire [3:0] deq_io_enq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] deq_io_enq_bits_prot; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] deq_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] deq_io_deq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] deq_io_deq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] deq_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] deq_io_deq_bits_burst; // @[Decoupled.scala 361:21]
  wire [3:0] deq_io_deq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] deq_io_deq_bits_prot; // @[Decoupled.scala 361:21]
  wire [29:0] deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  deq_metaReset; // @[Decoupled.scala 361:21]
  wire  deq_1_clock; // @[Decoupled.scala 361:21]
  wire  deq_1_reset; // @[Decoupled.scala 361:21]
  wire  deq_1_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  deq_1_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] deq_1_io_enq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] deq_1_io_enq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] deq_1_io_enq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] deq_1_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] deq_1_io_enq_bits_burst; // @[Decoupled.scala 361:21]
  wire [3:0] deq_1_io_enq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] deq_1_io_enq_bits_prot; // @[Decoupled.scala 361:21]
  wire  deq_1_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  deq_1_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [3:0] deq_1_io_deq_bits_id; // @[Decoupled.scala 361:21]
  wire [31:0] deq_1_io_deq_bits_addr; // @[Decoupled.scala 361:21]
  wire [7:0] deq_1_io_deq_bits_len; // @[Decoupled.scala 361:21]
  wire [2:0] deq_1_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [1:0] deq_1_io_deq_bits_burst; // @[Decoupled.scala 361:21]
  wire [3:0] deq_1_io_deq_bits_cache; // @[Decoupled.scala 361:21]
  wire [2:0] deq_1_io_deq_bits_prot; // @[Decoupled.scala 361:21]
  wire [29:0] deq_1_io_covSum; // @[Decoupled.scala 361:21]
  wire  deq_1_metaReset; // @[Decoupled.scala 361:21]
  wire  in_w_deq_clock; // @[Decoupled.scala 361:21]
  wire  in_w_deq_reset; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [63:0] in_w_deq_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] in_w_deq_io_enq_bits_strb; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_enq_bits_last; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [63:0] in_w_deq_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] in_w_deq_io_deq_bits_strb; // @[Decoupled.scala 361:21]
  wire  in_w_deq_io_deq_bits_last; // @[Decoupled.scala 361:21]
  wire [29:0] in_w_deq_io_covSum; // @[Decoupled.scala 361:21]
  wire  in_w_deq_metaReset; // @[Decoupled.scala 361:21]
  reg  busy; // @[Fragmenter.scala 60:29]
  reg [31:0] r_addr; // @[Fragmenter.scala 61:25]
  reg [7:0] r_len; // @[Fragmenter.scala 62:25]
  wire [7:0] irr_bits_len = deq_io_deq_bits_len; // @[Decoupled.scala 401:19 402:14]
  wire [7:0] len = busy ? r_len : irr_bits_len; // @[Fragmenter.scala 64:23]
  wire [31:0] irr_bits_addr = deq_io_deq_bits_addr; // @[Decoupled.scala 401:19 402:14]
  wire [31:0] addr = busy ? r_addr : irr_bits_addr; // @[Fragmenter.scala 65:23]
  wire [7:0] alignment = addr[10:3]; // @[Fragmenter.scala 69:29]
  wire [31:0] _support1_T = addr ^ 32'h2000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_1 = {1'b0,$signed(_support1_T)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_3 = $signed(_support1_T_1) & 33'sh86032000; // @[Parameters.scala 137:52]
  wire  _support1_T_4 = $signed(_support1_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  wire [32:0] _support1_T_6 = {1'b0,$signed(addr)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_8 = $signed(_support1_T_6) & 33'sh86012000; // @[Parameters.scala 137:52]
  wire  _support1_T_9 = $signed(_support1_T_8) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_10 = addr ^ 32'h10000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_11 = {1'b0,$signed(_support1_T_10)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_13 = $signed(_support1_T_11) & 33'sh86030000; // @[Parameters.scala 137:52]
  wire  _support1_T_14 = $signed(_support1_T_13) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_15 = addr ^ 32'h2000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_16 = {1'b0,$signed(_support1_T_15)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_18 = $signed(_support1_T_16) & 33'sh86030000; // @[Parameters.scala 137:52]
  wire  _support1_T_19 = $signed(_support1_T_18) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_20 = addr ^ 32'h4000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_21 = {1'b0,$signed(_support1_T_20)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_23 = $signed(_support1_T_21) & 33'sh84000000; // @[Parameters.scala 137:52]
  wire  _support1_T_24 = $signed(_support1_T_23) == 33'sh0; // @[Parameters.scala 137:67]
  wire [32:0] _support1_T_28 = $signed(_support1_T_21) & 33'sh86032000; // @[Parameters.scala 137:52]
  wire  _support1_T_29 = $signed(_support1_T_28) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_30 = addr ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_31 = {1'b0,$signed(_support1_T_30)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_33 = $signed(_support1_T_31) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  _support1_T_34 = $signed(_support1_T_33) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _support1_T_39 = _support1_T_9 | _support1_T_14 | _support1_T_19 | _support1_T_24 | _support1_T_29 |
    _support1_T_34; // @[Fragmenter.scala 76:100]
  wire [7:0] _support1_T_40 = _support1_T_4 ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [2:0] _support1_T_41 = _support1_T_39 ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [7:0] _GEN_44 = {{5'd0}, _support1_T_41}; // @[Mux.scala 27:73]
  wire [7:0] support1 = _support1_T_40 | _GEN_44; // @[Mux.scala 27:73]
  wire [7:0] _GEN_45 = {{1'd0}, len[7:1]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_1 = len | _GEN_45; // @[package.scala 253:43]
  wire [7:0] _GEN_46 = {{2'd0}, _fillLow_T_1[7:2]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_3 = _fillLow_T_1 | _GEN_46; // @[package.scala 253:43]
  wire [7:0] _GEN_47 = {{4'd0}, _fillLow_T_3[7:4]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_5 = _fillLow_T_3 | _GEN_47; // @[package.scala 253:43]
  wire [6:0] fillLow = _fillLow_T_5[7:1]; // @[Fragmenter.scala 85:37]
  wire [7:0] _wipeHigh_T = ~len; // @[Fragmenter.scala 86:32]
  wire [8:0] _wipeHigh_T_1 = {_wipeHigh_T, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_3 = _wipeHigh_T | _wipeHigh_T_1[7:0]; // @[package.scala 244:43]
  wire [9:0] _wipeHigh_T_4 = {_wipeHigh_T_3, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_6 = _wipeHigh_T_3 | _wipeHigh_T_4[7:0]; // @[package.scala 244:43]
  wire [11:0] _wipeHigh_T_7 = {_wipeHigh_T_6, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_9 = _wipeHigh_T_6 | _wipeHigh_T_7[7:0]; // @[package.scala 244:43]
  wire [7:0] wipeHigh = ~_wipeHigh_T_9; // @[Fragmenter.scala 86:24]
  wire [7:0] _GEN_48 = {{1'd0}, fillLow}; // @[Fragmenter.scala 87:32]
  wire [7:0] remain1 = _GEN_48 | wipeHigh; // @[Fragmenter.scala 87:32]
  wire [8:0] _align1_T = {alignment, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_2 = alignment | _align1_T[7:0]; // @[package.scala 244:43]
  wire [9:0] _align1_T_3 = {_align1_T_2, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_5 = _align1_T_2 | _align1_T_3[7:0]; // @[package.scala 244:43]
  wire [11:0] _align1_T_6 = {_align1_T_5, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_8 = _align1_T_5 | _align1_T_6[7:0]; // @[package.scala 244:43]
  wire [7:0] align1 = ~_align1_T_8; // @[Fragmenter.scala 88:24]
  wire [7:0] _maxSupported1_T = remain1 & align1; // @[Fragmenter.scala 89:37]
  wire [7:0] maxSupported1 = _maxSupported1_T & support1; // @[Fragmenter.scala 89:46]
  wire [1:0] irr_bits_burst = deq_io_deq_bits_burst; // @[Decoupled.scala 401:19 402:14]
  wire  fixed = irr_bits_burst == 2'h0; // @[Fragmenter.scala 92:34]
  wire [2:0] irr_bits_size = deq_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  wire  narrow = irr_bits_size != 3'h3; // @[Fragmenter.scala 93:34]
  wire  bad = fixed | narrow; // @[Fragmenter.scala 94:25]
  wire [7:0] beats1 = bad ? 8'h0 : maxSupported1; // @[Fragmenter.scala 97:25]
  wire [8:0] _beats_T = {beats1, 1'h0}; // @[package.scala 232:35]
  wire [8:0] _beats_T_1 = _beats_T | 9'h1; // @[package.scala 232:40]
  wire [8:0] _beats_T_2 = {1'h0,beats1}; // @[Cat.scala 31:58]
  wire [8:0] _beats_T_3 = ~_beats_T_2; // @[package.scala 232:53]
  wire [8:0] beats = _beats_T_1 & _beats_T_3; // @[package.scala 232:51]
  wire [15:0] _GEN_34 = {{7'd0}, beats}; // @[Fragmenter.scala 100:38]
  wire [15:0] _inc_addr_T = _GEN_34 << irr_bits_size; // @[Fragmenter.scala 100:38]
  wire [31:0] _GEN_49 = {{16'd0}, _inc_addr_T}; // @[Fragmenter.scala 100:29]
  wire [31:0] inc_addr = addr + _GEN_49; // @[Fragmenter.scala 100:29]
  wire [15:0] _wrapMask_T = {irr_bits_len,8'hff}; // @[Cat.scala 31:58]
  wire [22:0] _GEN_35 = {{7'd0}, _wrapMask_T}; // @[Bundles.scala 31:21]
  wire [22:0] _wrapMask_T_1 = _GEN_35 << irr_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] wrapMask = _wrapMask_T_1[22:8]; // @[Bundles.scala 31:30]
  wire [31:0] _GEN_50 = {{17'd0}, wrapMask}; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T = inc_addr & _GEN_50; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T_1 = ~irr_bits_addr; // @[Fragmenter.scala 104:49]
  wire [31:0] _mux_addr_T_2 = _mux_addr_T_1 | _GEN_50; // @[Fragmenter.scala 104:62]
  wire [31:0] _mux_addr_T_3 = ~_mux_addr_T_2; // @[Fragmenter.scala 104:47]
  wire [31:0] _mux_addr_T_4 = _mux_addr_T | _mux_addr_T_3; // @[Fragmenter.scala 104:45]
  wire  ar_last = beats1 == len; // @[Fragmenter.scala 110:27]
  wire [31:0] _out_bits_addr_T = ~addr; // @[Fragmenter.scala 122:28]
  wire [9:0] _out_bits_addr_T_2 = 10'h7 << irr_bits_size; // @[package.scala 234:77]
  wire [2:0] _out_bits_addr_T_4 = ~_out_bits_addr_T_2[2:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_52 = {{29'd0}, _out_bits_addr_T_4}; // @[Fragmenter.scala 122:34]
  wire [31:0] _out_bits_addr_T_5 = _out_bits_addr_T | _GEN_52; // @[Fragmenter.scala 122:34]
  wire  irr_valid = deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  wire  _T_2 = auto_out_ar_ready & irr_valid; // @[Decoupled.scala 50:35]
  wire [8:0] _GEN_53 = {{1'd0}, len}; // @[Fragmenter.scala 127:25]
  wire [8:0] _r_len_T_1 = _GEN_53 - beats; // @[Fragmenter.scala 127:25]
  wire [8:0] _GEN_4 = _T_2 ? _r_len_T_1 : {{1'd0}, r_len}; // @[Fragmenter.scala 124:27 127:18 62:25]
  reg  busy_1; // @[Fragmenter.scala 60:29]
  reg [31:0] r_addr_1; // @[Fragmenter.scala 61:25]
  reg [7:0] r_len_1; // @[Fragmenter.scala 62:25]
  wire [7:0] irr_1_bits_len = deq_1_io_deq_bits_len; // @[Decoupled.scala 401:19 402:14]
  wire [7:0] len_1 = busy_1 ? r_len_1 : irr_1_bits_len; // @[Fragmenter.scala 64:23]
  wire [31:0] irr_1_bits_addr = deq_1_io_deq_bits_addr; // @[Decoupled.scala 401:19 402:14]
  wire [31:0] addr_1 = busy_1 ? r_addr_1 : irr_1_bits_addr; // @[Fragmenter.scala 65:23]
  wire [7:0] alignment_1 = addr_1[10:3]; // @[Fragmenter.scala 69:29]
  wire [31:0] _support1_T_43 = addr_1 ^ 32'h2000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_44 = {1'b0,$signed(_support1_T_43)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_46 = $signed(_support1_T_44) & 33'sh86002000; // @[Parameters.scala 137:52]
  wire  _support1_T_47 = $signed(_support1_T_46) == 33'sh0; // @[Parameters.scala 137:67]
  wire [32:0] _support1_T_49 = {1'b0,$signed(addr_1)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_51 = $signed(_support1_T_49) & 33'sh82002000; // @[Parameters.scala 137:52]
  wire  _support1_T_52 = $signed(_support1_T_51) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_53 = addr_1 ^ 32'h2000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_54 = {1'b0,$signed(_support1_T_53)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_56 = $signed(_support1_T_54) & 33'sh86000000; // @[Parameters.scala 137:52]
  wire  _support1_T_57 = $signed(_support1_T_56) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_58 = addr_1 ^ 32'h4000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_59 = {1'b0,$signed(_support1_T_58)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_61 = $signed(_support1_T_59) & 33'sh84000000; // @[Parameters.scala 137:52]
  wire  _support1_T_62 = $signed(_support1_T_61) == 33'sh0; // @[Parameters.scala 137:67]
  wire [31:0] _support1_T_63 = addr_1 ^ 32'h80000000; // @[Parameters.scala 137:31]
  wire [32:0] _support1_T_64 = {1'b0,$signed(_support1_T_63)}; // @[Parameters.scala 137:49]
  wire [32:0] _support1_T_66 = $signed(_support1_T_64) & 33'sh80000000; // @[Parameters.scala 137:52]
  wire  _support1_T_67 = $signed(_support1_T_66) == 33'sh0; // @[Parameters.scala 137:67]
  wire  _support1_T_70 = _support1_T_52 | _support1_T_57 | _support1_T_62 | _support1_T_67; // @[Fragmenter.scala 76:100]
  wire [7:0] _support1_T_71 = _support1_T_47 ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [2:0] _support1_T_72 = _support1_T_70 ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [7:0] _GEN_54 = {{5'd0}, _support1_T_72}; // @[Mux.scala 27:73]
  wire [7:0] support1_1 = _support1_T_71 | _GEN_54; // @[Mux.scala 27:73]
  wire [7:0] _GEN_55 = {{1'd0}, len_1[7:1]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_8 = len_1 | _GEN_55; // @[package.scala 253:43]
  wire [7:0] _GEN_56 = {{2'd0}, _fillLow_T_8[7:2]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_10 = _fillLow_T_8 | _GEN_56; // @[package.scala 253:43]
  wire [7:0] _GEN_57 = {{4'd0}, _fillLow_T_10[7:4]}; // @[package.scala 253:43]
  wire [7:0] _fillLow_T_12 = _fillLow_T_10 | _GEN_57; // @[package.scala 253:43]
  wire [6:0] fillLow_1 = _fillLow_T_12[7:1]; // @[Fragmenter.scala 85:37]
  wire [7:0] _wipeHigh_T_11 = ~len_1; // @[Fragmenter.scala 86:32]
  wire [8:0] _wipeHigh_T_12 = {_wipeHigh_T_11, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_14 = _wipeHigh_T_11 | _wipeHigh_T_12[7:0]; // @[package.scala 244:43]
  wire [9:0] _wipeHigh_T_15 = {_wipeHigh_T_14, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_17 = _wipeHigh_T_14 | _wipeHigh_T_15[7:0]; // @[package.scala 244:43]
  wire [11:0] _wipeHigh_T_18 = {_wipeHigh_T_17, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _wipeHigh_T_20 = _wipeHigh_T_17 | _wipeHigh_T_18[7:0]; // @[package.scala 244:43]
  wire [7:0] wipeHigh_1 = ~_wipeHigh_T_20; // @[Fragmenter.scala 86:24]
  wire [7:0] _GEN_58 = {{1'd0}, fillLow_1}; // @[Fragmenter.scala 87:32]
  wire [7:0] remain1_1 = _GEN_58 | wipeHigh_1; // @[Fragmenter.scala 87:32]
  wire [8:0] _align1_T_10 = {alignment_1, 1'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_12 = alignment_1 | _align1_T_10[7:0]; // @[package.scala 244:43]
  wire [9:0] _align1_T_13 = {_align1_T_12, 2'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_15 = _align1_T_12 | _align1_T_13[7:0]; // @[package.scala 244:43]
  wire [11:0] _align1_T_16 = {_align1_T_15, 4'h0}; // @[package.scala 244:48]
  wire [7:0] _align1_T_18 = _align1_T_15 | _align1_T_16[7:0]; // @[package.scala 244:43]
  wire [7:0] align1_1 = ~_align1_T_18; // @[Fragmenter.scala 88:24]
  wire [7:0] _maxSupported1_T_1 = remain1_1 & align1_1; // @[Fragmenter.scala 89:37]
  wire [7:0] maxSupported1_1 = _maxSupported1_T_1 & support1_1; // @[Fragmenter.scala 89:46]
  wire [1:0] irr_1_bits_burst = deq_1_io_deq_bits_burst; // @[Decoupled.scala 401:19 402:14]
  wire  fixed_1 = irr_1_bits_burst == 2'h0; // @[Fragmenter.scala 92:34]
  wire [2:0] irr_1_bits_size = deq_1_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  wire  narrow_1 = irr_1_bits_size != 3'h3; // @[Fragmenter.scala 93:34]
  wire  bad_1 = fixed_1 | narrow_1; // @[Fragmenter.scala 94:25]
  wire [7:0] beats1_1 = bad_1 ? 8'h0 : maxSupported1_1; // @[Fragmenter.scala 97:25]
  wire [8:0] _beats_T_4 = {beats1_1, 1'h0}; // @[package.scala 232:35]
  wire [8:0] _beats_T_5 = _beats_T_4 | 9'h1; // @[package.scala 232:40]
  wire [8:0] _beats_T_6 = {1'h0,beats1_1}; // @[Cat.scala 31:58]
  wire [8:0] _beats_T_7 = ~_beats_T_6; // @[package.scala 232:53]
  wire [8:0] w_beats = _beats_T_5 & _beats_T_7; // @[package.scala 232:51]
  wire [15:0] _GEN_70 = {{7'd0}, w_beats}; // @[Fragmenter.scala 100:38]
  wire [15:0] _inc_addr_T_2 = _GEN_70 << irr_1_bits_size; // @[Fragmenter.scala 100:38]
  wire [31:0] _GEN_59 = {{16'd0}, _inc_addr_T_2}; // @[Fragmenter.scala 100:29]
  wire [31:0] inc_addr_1 = addr_1 + _GEN_59; // @[Fragmenter.scala 100:29]
  wire [15:0] _wrapMask_T_2 = {irr_1_bits_len,8'hff}; // @[Cat.scala 31:58]
  wire [22:0] _GEN_71 = {{7'd0}, _wrapMask_T_2}; // @[Bundles.scala 31:21]
  wire [22:0] _wrapMask_T_3 = _GEN_71 << irr_1_bits_size; // @[Bundles.scala 31:21]
  wire [14:0] wrapMask_1 = _wrapMask_T_3[22:8]; // @[Bundles.scala 31:30]
  wire [31:0] _GEN_60 = {{17'd0}, wrapMask_1}; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T_5 = inc_addr_1 & _GEN_60; // @[Fragmenter.scala 104:33]
  wire [31:0] _mux_addr_T_6 = ~irr_1_bits_addr; // @[Fragmenter.scala 104:49]
  wire [31:0] _mux_addr_T_7 = _mux_addr_T_6 | _GEN_60; // @[Fragmenter.scala 104:62]
  wire [31:0] _mux_addr_T_8 = ~_mux_addr_T_7; // @[Fragmenter.scala 104:47]
  wire [31:0] _mux_addr_T_9 = _mux_addr_T_5 | _mux_addr_T_8; // @[Fragmenter.scala 104:45]
  wire  aw_last = beats1_1 == len_1; // @[Fragmenter.scala 110:27]
  reg [8:0] w_counter; // @[Fragmenter.scala 164:30]
  wire  w_idle = w_counter == 9'h0; // @[Fragmenter.scala 165:30]
  reg  wbeats_latched; // @[Fragmenter.scala 150:35]
  wire  _in_aw_ready_T = w_idle | wbeats_latched; // @[Fragmenter.scala 158:52]
  wire  in_aw_ready = auto_out_aw_ready & (w_idle | wbeats_latched); // @[Fragmenter.scala 158:35]
  wire [31:0] _out_bits_addr_T_7 = ~addr_1; // @[Fragmenter.scala 122:28]
  wire [9:0] _out_bits_addr_T_9 = 10'h7 << irr_1_bits_size; // @[package.scala 234:77]
  wire [2:0] _out_bits_addr_T_11 = ~_out_bits_addr_T_9[2:0]; // @[package.scala 234:46]
  wire [31:0] _GEN_62 = {{29'd0}, _out_bits_addr_T_11}; // @[Fragmenter.scala 122:34]
  wire [31:0] _out_bits_addr_T_12 = _out_bits_addr_T_7 | _GEN_62; // @[Fragmenter.scala 122:34]
  wire  irr_1_valid = deq_1_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  wire  _T_5 = in_aw_ready & irr_1_valid; // @[Decoupled.scala 50:35]
  wire [8:0] _GEN_63 = {{1'd0}, len_1}; // @[Fragmenter.scala 127:25]
  wire [8:0] _r_len_T_3 = _GEN_63 - w_beats; // @[Fragmenter.scala 127:25]
  wire [8:0] _GEN_9 = _T_5 ? _r_len_T_3 : {{1'd0}, r_len_1}; // @[Fragmenter.scala 124:27 127:18 62:25]
  wire  wbeats_valid = irr_1_valid & ~wbeats_latched; // @[Fragmenter.scala 159:35]
  wire  _GEN_10 = wbeats_valid & w_idle | wbeats_latched; // @[Fragmenter.scala 150:35 153:{43,60}]
  wire  bundleOut_0_aw_valid = irr_1_valid & _in_aw_ready_T; // @[Fragmenter.scala 157:35]
  wire  _T_7 = auto_out_aw_ready & bundleOut_0_aw_valid; // @[Decoupled.scala 50:35]
  wire [8:0] _w_todo_T = wbeats_valid ? w_beats : 9'h0; // @[Fragmenter.scala 166:35]
  wire [8:0] w_todo = w_idle ? _w_todo_T : w_counter; // @[Fragmenter.scala 166:23]
  wire  w_last = w_todo == 9'h1; // @[Fragmenter.scala 167:27]
  wire  in_w_valid = in_w_deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  wire  _bundleOut_0_w_valid_T_1 = ~w_idle | wbeats_valid; // @[Fragmenter.scala 173:51]
  wire  bundleOut_0_w_valid = in_w_valid & (~w_idle | wbeats_valid); // @[Fragmenter.scala 173:33]
  wire  _w_counter_T = auto_out_w_ready & bundleOut_0_w_valid; // @[Decoupled.scala 50:35]
  wire [8:0] _GEN_64 = {{8'd0}, _w_counter_T}; // @[Fragmenter.scala 168:27]
  wire [8:0] _w_counter_T_2 = w_todo - _GEN_64; // @[Fragmenter.scala 168:27]
  wire  _T_13 = ~reset; // @[Fragmenter.scala 169:14]
  wire  in_w_bits_last = in_w_deq_io_deq_bits_last; // @[Decoupled.scala 401:19 402:14]
  wire  bundleOut_0_b_ready = auto_in_b_ready | ~auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 189:33]
  reg [1:0] error_0; // @[Fragmenter.scala 192:26]
  reg [1:0] error_1; // @[Fragmenter.scala 192:26]
  reg [1:0] error_2; // @[Fragmenter.scala 192:26]
  reg [1:0] error_3; // @[Fragmenter.scala 192:26]
  reg [1:0] error_4; // @[Fragmenter.scala 192:26]
  reg [1:0] error_5; // @[Fragmenter.scala 192:26]
  reg [1:0] error_6; // @[Fragmenter.scala 192:26]
  reg [1:0] error_7; // @[Fragmenter.scala 192:26]
  reg [1:0] error_8; // @[Fragmenter.scala 192:26]
  reg [1:0] error_9; // @[Fragmenter.scala 192:26]
  reg [1:0] error_10; // @[Fragmenter.scala 192:26]
  reg [1:0] error_11; // @[Fragmenter.scala 192:26]
  reg [1:0] error_12; // @[Fragmenter.scala 192:26]
  reg [1:0] error_13; // @[Fragmenter.scala 192:26]
  reg [1:0] error_14; // @[Fragmenter.scala 192:26]
  reg [1:0] error_15; // @[Fragmenter.scala 192:26]
  wire [1:0] _GEN_13 = 4'h1 == auto_out_b_bits_id ? error_1 : error_0; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_14 = 4'h2 == auto_out_b_bits_id ? error_2 : _GEN_13; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_15 = 4'h3 == auto_out_b_bits_id ? error_3 : _GEN_14; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_16 = 4'h4 == auto_out_b_bits_id ? error_4 : _GEN_15; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_17 = 4'h5 == auto_out_b_bits_id ? error_5 : _GEN_16; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_18 = 4'h6 == auto_out_b_bits_id ? error_6 : _GEN_17; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_19 = 4'h7 == auto_out_b_bits_id ? error_7 : _GEN_18; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_20 = 4'h8 == auto_out_b_bits_id ? error_8 : _GEN_19; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_21 = 4'h9 == auto_out_b_bits_id ? error_9 : _GEN_20; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_22 = 4'ha == auto_out_b_bits_id ? error_10 : _GEN_21; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_23 = 4'hb == auto_out_b_bits_id ? error_11 : _GEN_22; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_24 = 4'hc == auto_out_b_bits_id ? error_12 : _GEN_23; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_25 = 4'hd == auto_out_b_bits_id ? error_13 : _GEN_24; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_26 = 4'he == auto_out_b_bits_id ? error_14 : _GEN_25; // @[Fragmenter.scala 193:{41,41}]
  wire [1:0] _GEN_27 = 4'hf == auto_out_b_bits_id ? error_15 : _GEN_26; // @[Fragmenter.scala 193:{41,41}]
  wire [15:0] _T_22 = 16'h1 << auto_out_b_bits_id; // @[OneHot.scala 64:12]
  wire  _T_40 = bundleOut_0_b_ready & auto_out_b_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _error_0_T = error_0 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_1_T = error_1 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_2_T = error_2 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_3_T = error_3 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_4_T = error_4 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_5_T = error_5 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_6_T = error_6 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_7_T = error_7 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_8_T = error_8 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_9_T = error_9 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_10_T = error_10 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_11_T = error_11 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_12_T = error_12 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_13_T = error_13 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_14_T = error_14 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  wire [1:0] _error_15_T = error_15 | auto_out_b_bits_resp; // @[Fragmenter.scala 195:70]
  reg [6:0] AXI4Fragmenter_1_covState; // @[Register tracking AXI4Fragmenter_1 state]
  reg  AXI4Fragmenter_1_covMap [0:127]; // @[Coverage map for AXI4Fragmenter_1]
  wire  AXI4Fragmenter_1_covMap_read_en; // @[Coverage map for AXI4Fragmenter_1]
  wire [6:0] AXI4Fragmenter_1_covMap_read_addr; // @[Coverage map for AXI4Fragmenter_1]
  wire  AXI4Fragmenter_1_covMap_read_data; // @[Coverage map for AXI4Fragmenter_1]
  wire  AXI4Fragmenter_1_covMap_write_data; // @[Coverage map for AXI4Fragmenter_1]
  wire [6:0] AXI4Fragmenter_1_covMap_write_addr; // @[Coverage map for AXI4Fragmenter_1]
  wire  AXI4Fragmenter_1_covMap_write_mask; // @[Coverage map for AXI4Fragmenter_1]
  wire  AXI4Fragmenter_1_covMap_write_en; // @[Coverage map for AXI4Fragmenter_1]
  reg [29:0] AXI4Fragmenter_1_covSum; // @[Sum of coverage map]
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  busy_shl;
  wire [6:0] busy_pad;
  wire [1:0] wbeats_latched_shl;
  wire [6:0] wbeats_latched_pad;
  wire [2:0] busy_1_shl;
  wire [6:0] busy_1_pad;
  wire [3:0] mux_cond_0_shl;
  wire [6:0] mux_cond_0_pad;
  wire [4:0] mux_cond_1_shl;
  wire [6:0] mux_cond_1_pad;
  wire [5:0] mux_cond_2_shl;
  wire [6:0] mux_cond_2_pad;
  wire [6:0] mux_cond_3_shl;
  wire [6:0] mux_cond_3_pad;
  wire [6:0] AXI4Fragmenter_1_xor4;
  wire [6:0] AXI4Fragmenter_1_xor1;
  wire [6:0] AXI4Fragmenter_1_xor5;
  wire [6:0] AXI4Fragmenter_1_xor6;
  wire [6:0] AXI4Fragmenter_1_xor2;
  wire [6:0] AXI4Fragmenter_1_xor0;
  wire [29:0] deq_sum;
  wire [29:0] deq_1_sum;
  wire [29:0] in_w_deq_sum;
  Queue_28 deq ( // @[Decoupled.scala 361:21]
    .clock(deq_clock),
    .reset(deq_reset),
    .io_enq_ready(deq_io_enq_ready),
    .io_enq_valid(deq_io_enq_valid),
    .io_enq_bits_id(deq_io_enq_bits_id),
    .io_enq_bits_addr(deq_io_enq_bits_addr),
    .io_enq_bits_len(deq_io_enq_bits_len),
    .io_enq_bits_size(deq_io_enq_bits_size),
    .io_enq_bits_burst(deq_io_enq_bits_burst),
    .io_enq_bits_cache(deq_io_enq_bits_cache),
    .io_enq_bits_prot(deq_io_enq_bits_prot),
    .io_deq_ready(deq_io_deq_ready),
    .io_deq_valid(deq_io_deq_valid),
    .io_deq_bits_id(deq_io_deq_bits_id),
    .io_deq_bits_addr(deq_io_deq_bits_addr),
    .io_deq_bits_len(deq_io_deq_bits_len),
    .io_deq_bits_size(deq_io_deq_bits_size),
    .io_deq_bits_burst(deq_io_deq_bits_burst),
    .io_deq_bits_cache(deq_io_deq_bits_cache),
    .io_deq_bits_prot(deq_io_deq_bits_prot),
    .io_covSum(deq_io_covSum),
    .metaReset(deq_metaReset)
  );
  Queue_28 deq_1 ( // @[Decoupled.scala 361:21]
    .clock(deq_1_clock),
    .reset(deq_1_reset),
    .io_enq_ready(deq_1_io_enq_ready),
    .io_enq_valid(deq_1_io_enq_valid),
    .io_enq_bits_id(deq_1_io_enq_bits_id),
    .io_enq_bits_addr(deq_1_io_enq_bits_addr),
    .io_enq_bits_len(deq_1_io_enq_bits_len),
    .io_enq_bits_size(deq_1_io_enq_bits_size),
    .io_enq_bits_burst(deq_1_io_enq_bits_burst),
    .io_enq_bits_cache(deq_1_io_enq_bits_cache),
    .io_enq_bits_prot(deq_1_io_enq_bits_prot),
    .io_deq_ready(deq_1_io_deq_ready),
    .io_deq_valid(deq_1_io_deq_valid),
    .io_deq_bits_id(deq_1_io_deq_bits_id),
    .io_deq_bits_addr(deq_1_io_deq_bits_addr),
    .io_deq_bits_len(deq_1_io_deq_bits_len),
    .io_deq_bits_size(deq_1_io_deq_bits_size),
    .io_deq_bits_burst(deq_1_io_deq_bits_burst),
    .io_deq_bits_cache(deq_1_io_deq_bits_cache),
    .io_deq_bits_prot(deq_1_io_deq_bits_prot),
    .io_covSum(deq_1_io_covSum),
    .metaReset(deq_1_metaReset)
  );
  Queue_12 in_w_deq ( // @[Decoupled.scala 361:21]
    .clock(in_w_deq_clock),
    .reset(in_w_deq_reset),
    .io_enq_ready(in_w_deq_io_enq_ready),
    .io_enq_valid(in_w_deq_io_enq_valid),
    .io_enq_bits_data(in_w_deq_io_enq_bits_data),
    .io_enq_bits_strb(in_w_deq_io_enq_bits_strb),
    .io_enq_bits_last(in_w_deq_io_enq_bits_last),
    .io_deq_ready(in_w_deq_io_deq_ready),
    .io_deq_valid(in_w_deq_io_deq_valid),
    .io_deq_bits_data(in_w_deq_io_deq_bits_data),
    .io_deq_bits_strb(in_w_deq_io_deq_bits_strb),
    .io_deq_bits_last(in_w_deq_io_deq_bits_last),
    .io_covSum(in_w_deq_io_covSum),
    .metaReset(in_w_deq_metaReset)
  );
  assign auto_in_aw_ready = deq_1_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_w_ready = in_w_deq_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_b_valid = auto_out_b_valid & auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 188:33]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp | _GEN_27; // @[Fragmenter.scala 193:41]
  assign auto_in_ar_ready = deq_io_enq_ready; // @[Nodes.scala 1210:84 Decoupled.scala 365:17]
  assign auto_in_r_valid = auto_out_r_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last & auto_out_r_bits_echo_real_last; // @[Fragmenter.scala 183:41]
  assign auto_out_aw_valid = irr_1_valid & _in_aw_ready_T; // @[Fragmenter.scala 157:35]
  assign auto_out_aw_bits_id = deq_1_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_addr = ~_out_bits_addr_T_12; // @[Fragmenter.scala 122:26]
  assign auto_out_aw_bits_len = bad_1 ? 8'h0 : maxSupported1_1; // @[Fragmenter.scala 97:25]
  assign auto_out_aw_bits_size = deq_1_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_cache = deq_1_io_deq_bits_cache; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_prot = deq_1_io_deq_bits_prot; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_aw_bits_echo_real_last = beats1_1 == len_1; // @[Fragmenter.scala 110:27]
  assign auto_out_w_valid = in_w_valid & (~w_idle | wbeats_valid); // @[Fragmenter.scala 173:33]
  assign auto_out_w_bits_data = in_w_deq_io_deq_bits_data; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_w_bits_strb = in_w_deq_io_deq_bits_strb; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_w_bits_last = w_todo == 9'h1; // @[Fragmenter.scala 167:27]
  assign auto_out_b_ready = auto_in_b_ready | ~auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 189:33]
  assign auto_out_ar_valid = deq_io_deq_valid; // @[Decoupled.scala 401:19 403:15]
  assign auto_out_ar_bits_id = deq_io_deq_bits_id; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_addr = ~_out_bits_addr_T_5; // @[Fragmenter.scala 122:26]
  assign auto_out_ar_bits_len = bad ? 8'h0 : maxSupported1; // @[Fragmenter.scala 97:25]
  assign auto_out_ar_bits_size = deq_io_deq_bits_size; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_cache = deq_io_deq_bits_cache; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_prot = deq_io_deq_bits_prot; // @[Decoupled.scala 401:19 402:14]
  assign auto_out_ar_bits_echo_real_last = beats1 == len; // @[Fragmenter.scala 110:27]
  assign auto_out_r_ready = auto_in_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_clock = clock;
  assign deq_reset = reset;
  assign deq_io_enq_valid = auto_in_ar_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_id = auto_in_ar_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_len = auto_in_ar_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_size = auto_in_ar_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_burst = auto_in_ar_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_cache = auto_in_ar_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_enq_bits_prot = auto_in_ar_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_io_deq_ready = auto_out_ar_ready & ar_last; // @[Fragmenter.scala 111:30]
  assign deq_1_clock = clock;
  assign deq_1_reset = reset;
  assign deq_1_io_enq_valid = auto_in_aw_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_id = auto_in_aw_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_len = auto_in_aw_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_size = auto_in_aw_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_burst = auto_in_aw_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_cache = auto_in_aw_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_enq_bits_prot = auto_in_aw_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign deq_1_io_deq_ready = in_aw_ready & aw_last; // @[Fragmenter.scala 111:30]
  assign in_w_deq_clock = clock;
  assign in_w_deq_reset = reset;
  assign in_w_deq_io_enq_valid = auto_in_w_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_w_deq_io_enq_bits_data = auto_in_w_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_w_deq_io_enq_bits_strb = auto_in_w_bits_strb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_w_deq_io_enq_bits_last = auto_in_w_bits_last; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign in_w_deq_io_deq_ready = auto_out_w_ready & _bundleOut_0_w_valid_T_1; // @[Fragmenter.scala 174:33]
  assign AXI4Fragmenter_1_covMap_read_en = 1'h1;
  assign AXI4Fragmenter_1_covMap_read_addr = AXI4Fragmenter_1_covState;
  assign AXI4Fragmenter_1_covMap_read_data = AXI4Fragmenter_1_covMap[AXI4Fragmenter_1_covMap_read_addr]; // @[Coverage map for AXI4Fragmenter_1]
  assign AXI4Fragmenter_1_covMap_write_data = 1'h1;
  assign AXI4Fragmenter_1_covMap_write_addr = AXI4Fragmenter_1_covState;
  assign AXI4Fragmenter_1_covMap_write_mask = 1'h1;
  assign AXI4Fragmenter_1_covMap_write_en = ~metaReset;
  assign mux_cond_0 = _support1_T_47;
  assign mux_cond_1 = _support1_T_4;
  assign mux_cond_2 = _support1_T_39;
  assign mux_cond_3 = _support1_T_70;
  assign busy_shl = busy;
  assign busy_pad = {6'h0,busy_shl};
  assign wbeats_latched_shl = {wbeats_latched, 1'h0};
  assign wbeats_latched_pad = {5'h0,wbeats_latched_shl};
  assign busy_1_shl = {busy_1, 2'h0};
  assign busy_1_pad = {4'h0,busy_1_shl};
  assign mux_cond_0_shl = {mux_cond_0, 3'h0};
  assign mux_cond_0_pad = {3'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 4'h0};
  assign mux_cond_1_pad = {2'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 5'h0};
  assign mux_cond_2_pad = {1'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 6'h0};
  assign mux_cond_3_pad = mux_cond_3_shl;
  assign AXI4Fragmenter_1_xor4 = wbeats_latched_pad ^ busy_1_pad;
  assign AXI4Fragmenter_1_xor1 = busy_pad ^ AXI4Fragmenter_1_xor4;
  assign AXI4Fragmenter_1_xor5 = mux_cond_0_pad ^ mux_cond_1_pad;
  assign AXI4Fragmenter_1_xor6 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign AXI4Fragmenter_1_xor2 = AXI4Fragmenter_1_xor5 ^ AXI4Fragmenter_1_xor6;
  assign AXI4Fragmenter_1_xor0 = AXI4Fragmenter_1_xor1 ^ AXI4Fragmenter_1_xor2;
  assign deq_sum = AXI4Fragmenter_1_covSum + deq_io_covSum;
  assign deq_1_sum = deq_sum + deq_1_io_covSum;
  assign in_w_deq_sum = deq_1_sum + in_w_deq_io_covSum;
  assign io_covSum = in_w_deq_sum;
  assign deq_metaReset = metaReset;
  assign deq_1_metaReset = metaReset;
  assign in_w_deq_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 60:29]
      busy <= 1'h0; // @[Fragmenter.scala 60:29]
    end else if (_T_2) begin
      busy <= ~ar_last;
    end
    if (_T_2) begin // @[Fragmenter.scala 124:27]
      if (fixed) begin
        r_addr <= irr_bits_addr;
      end else if (irr_bits_burst == 2'h2) begin
        r_addr <= _mux_addr_T_4;
      end else begin
        r_addr <= inc_addr;
      end
    end
    r_len <= _GEN_4[7:0];
    if (reset) begin // @[Fragmenter.scala 60:29]
      busy_1 <= 1'h0; // @[Fragmenter.scala 60:29]
    end else if (_T_5) begin
      busy_1 <= ~aw_last;
    end
    if (_T_5) begin // @[Fragmenter.scala 124:27]
      if (fixed_1) begin
        r_addr_1 <= irr_1_bits_addr;
      end else if (irr_1_bits_burst == 2'h2) begin
        r_addr_1 <= _mux_addr_T_9;
      end else begin
        r_addr_1 <= inc_addr_1;
      end
    end
    r_len_1 <= _GEN_9[7:0];
    if (reset) begin // @[Fragmenter.scala 164:30]
      w_counter <= 9'h0; // @[Fragmenter.scala 164:30]
    end else begin
      w_counter <= _w_counter_T_2; // @[Fragmenter.scala 168:17]
    end
    if (reset) begin // @[Fragmenter.scala 150:35]
      wbeats_latched <= 1'h0; // @[Fragmenter.scala 150:35]
    end else if (_T_7) begin
      wbeats_latched <= 1'h0;
    end else begin
      wbeats_latched <= _GEN_10;
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_0 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[0] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_0 <= 2'h0;
      end else begin
        error_0 <= _error_0_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_1 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[1] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_1 <= 2'h0;
      end else begin
        error_1 <= _error_1_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_2 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[2] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_2 <= 2'h0;
      end else begin
        error_2 <= _error_2_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_3 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[3] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_3 <= 2'h0;
      end else begin
        error_3 <= _error_3_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_4 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[4] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_4 <= 2'h0;
      end else begin
        error_4 <= _error_4_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_5 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[5] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_5 <= 2'h0;
      end else begin
        error_5 <= _error_5_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_6 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[6] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_6 <= 2'h0;
      end else begin
        error_6 <= _error_6_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_7 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[7] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_7 <= 2'h0;
      end else begin
        error_7 <= _error_7_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_8 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[8] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_8 <= 2'h0;
      end else begin
        error_8 <= _error_8_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_9 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[9] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_9 <= 2'h0;
      end else begin
        error_9 <= _error_9_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_10 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[10] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_10 <= 2'h0;
      end else begin
        error_10 <= _error_10_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_11 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[11] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_11 <= 2'h0;
      end else begin
        error_11 <= _error_11_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_12 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[12] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_12 <= 2'h0;
      end else begin
        error_12 <= _error_12_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_13 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[13] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_13 <= 2'h0;
      end else begin
        error_13 <= _error_13_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_14 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[14] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_14 <= 2'h0;
      end else begin
        error_14 <= _error_14_T;
      end
    end
    if (reset) begin // @[Fragmenter.scala 192:26]
      error_15 <= 2'h0; // @[Fragmenter.scala 192:26]
    end else if (_T_22[15] & _T_40) begin
      if (auto_out_b_bits_echo_real_last) begin
        error_15 <= 2'h0;
      end else begin
        error_15 <= _error_15_T;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_w_counter_T | w_todo != 9'h0) & ~reset) begin
          $fatal; // @[Fragmenter.scala 169:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~_w_counter_T | w_todo != 9'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:169 assert (!out.w.fire() || w_todo =/= UInt(0)) // underflow impossible\n"
            ); // @[Fragmenter.scala 169:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~bundleOut_0_w_valid | ~in_w_bits_last | w_last) & _T_13) begin
          $fatal; // @[Fragmenter.scala 178:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(~bundleOut_0_w_valid | ~in_w_bits_last | w_last)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:178 assert (!out.w.valid || !in_w.bits.last || w_last)\n"); // @[Fragmenter.scala 178:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    AXI4Fragmenter_1_covState <= AXI4Fragmenter_1_xor0;
    if (AXI4Fragmenter_1_covMap_write_en & AXI4Fragmenter_1_covMap_write_mask) begin
      AXI4Fragmenter_1_covMap[AXI4Fragmenter_1_covMap_write_addr] <= AXI4Fragmenter_1_covMap_write_data; // @[Coverage map for AXI4Fragmenter_1]
    end
    if (!(AXI4Fragmenter_1_covMap_read_data | metaReset)) begin
      AXI4Fragmenter_1_covSum <= AXI4Fragmenter_1_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    AXI4Fragmenter_1_covMap[initvar] = 0; //_25[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_len = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  busy_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_addr_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  r_len_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  w_counter = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  wbeats_latched = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  error_0 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  error_1 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  error_2 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  error_3 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  error_4 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  error_5 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  error_6 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  error_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  error_8 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  error_9 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  error_10 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  error_11 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  error_12 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  error_13 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  error_14 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  error_15 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  AXI4Fragmenter_1_covState = 0; //_24[6:0];
  _RAND_26 = {1{`RANDOM}};
  AXI4Fragmenter_1_covSum = 0; //_26[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CVA6Tile(
  input         clock,
  input         reset,
  input         auto_int_local_in_3_0,
  input         auto_int_local_in_2_0,
  input         auto_int_local_in_1_0,
  input         auto_int_local_in_1_1,
  input         auto_hartid_in,
  input         auto_tl_other_masters_out_a_ready,
  output        auto_tl_other_masters_out_a_valid,
  output [2:0]  auto_tl_other_masters_out_a_bits_opcode,
  output [2:0]  auto_tl_other_masters_out_a_bits_param,
  output [3:0]  auto_tl_other_masters_out_a_bits_size,
  output [5:0]  auto_tl_other_masters_out_a_bits_source,
  output [31:0] auto_tl_other_masters_out_a_bits_address,
  output        auto_tl_other_masters_out_a_bits_user_amba_prot_bufferable,
  output        auto_tl_other_masters_out_a_bits_user_amba_prot_modifiable,
  output        auto_tl_other_masters_out_a_bits_user_amba_prot_readalloc,
  output        auto_tl_other_masters_out_a_bits_user_amba_prot_writealloc,
  output        auto_tl_other_masters_out_a_bits_user_amba_prot_privileged,
  output        auto_tl_other_masters_out_a_bits_user_amba_prot_secure,
  output        auto_tl_other_masters_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_tl_other_masters_out_a_bits_mask,
  output [63:0] auto_tl_other_masters_out_a_bits_data,
  output        auto_tl_other_masters_out_d_ready,
  input         auto_tl_other_masters_out_d_valid,
  input  [2:0]  auto_tl_other_masters_out_d_bits_opcode,
  input  [3:0]  auto_tl_other_masters_out_d_bits_size,
  input  [5:0]  auto_tl_other_masters_out_d_bits_source,
  input         auto_tl_other_masters_out_d_bits_denied,
  input  [63:0] auto_tl_other_masters_out_d_bits_data,
  input         auto_tl_other_masters_out_d_bits_corrupt,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  tlMasterXbar_auto_in_a_ready;
  wire  tlMasterXbar_auto_in_a_valid;
  wire [2:0] tlMasterXbar_auto_in_a_bits_opcode;
  wire [2:0] tlMasterXbar_auto_in_a_bits_param;
  wire [3:0] tlMasterXbar_auto_in_a_bits_size;
  wire [5:0] tlMasterXbar_auto_in_a_bits_source;
  wire [31:0] tlMasterXbar_auto_in_a_bits_address;
  wire  tlMasterXbar_auto_in_a_bits_user_amba_prot_bufferable;
  wire  tlMasterXbar_auto_in_a_bits_user_amba_prot_modifiable;
  wire  tlMasterXbar_auto_in_a_bits_user_amba_prot_readalloc;
  wire  tlMasterXbar_auto_in_a_bits_user_amba_prot_writealloc;
  wire  tlMasterXbar_auto_in_a_bits_user_amba_prot_privileged;
  wire  tlMasterXbar_auto_in_a_bits_user_amba_prot_secure;
  wire  tlMasterXbar_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] tlMasterXbar_auto_in_a_bits_mask;
  wire [63:0] tlMasterXbar_auto_in_a_bits_data;
  wire  tlMasterXbar_auto_in_d_ready;
  wire  tlMasterXbar_auto_in_d_valid;
  wire [2:0] tlMasterXbar_auto_in_d_bits_opcode;
  wire [3:0] tlMasterXbar_auto_in_d_bits_size;
  wire [5:0] tlMasterXbar_auto_in_d_bits_source;
  wire  tlMasterXbar_auto_in_d_bits_denied;
  wire [63:0] tlMasterXbar_auto_in_d_bits_data;
  wire  tlMasterXbar_auto_in_d_bits_corrupt;
  wire  tlMasterXbar_auto_out_a_ready;
  wire  tlMasterXbar_auto_out_a_valid;
  wire [2:0] tlMasterXbar_auto_out_a_bits_opcode;
  wire [2:0] tlMasterXbar_auto_out_a_bits_param;
  wire [3:0] tlMasterXbar_auto_out_a_bits_size;
  wire [5:0] tlMasterXbar_auto_out_a_bits_source;
  wire [31:0] tlMasterXbar_auto_out_a_bits_address;
  wire  tlMasterXbar_auto_out_a_bits_user_amba_prot_bufferable;
  wire  tlMasterXbar_auto_out_a_bits_user_amba_prot_modifiable;
  wire  tlMasterXbar_auto_out_a_bits_user_amba_prot_readalloc;
  wire  tlMasterXbar_auto_out_a_bits_user_amba_prot_writealloc;
  wire  tlMasterXbar_auto_out_a_bits_user_amba_prot_privileged;
  wire  tlMasterXbar_auto_out_a_bits_user_amba_prot_secure;
  wire  tlMasterXbar_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] tlMasterXbar_auto_out_a_bits_mask;
  wire [63:0] tlMasterXbar_auto_out_a_bits_data;
  wire  tlMasterXbar_auto_out_d_ready;
  wire  tlMasterXbar_auto_out_d_valid;
  wire [2:0] tlMasterXbar_auto_out_d_bits_opcode;
  wire [3:0] tlMasterXbar_auto_out_d_bits_size;
  wire [5:0] tlMasterXbar_auto_out_d_bits_source;
  wire  tlMasterXbar_auto_out_d_bits_denied;
  wire [63:0] tlMasterXbar_auto_out_d_bits_data;
  wire  tlMasterXbar_auto_out_d_bits_corrupt;
  wire  intXbar_auto_int_in_3_0; // @[BaseTile.scala 212:37]
  wire  intXbar_auto_int_in_2_0; // @[BaseTile.scala 212:37]
  wire  intXbar_auto_int_in_1_0; // @[BaseTile.scala 212:37]
  wire  intXbar_auto_int_in_1_1; // @[BaseTile.scala 212:37]
  wire  intXbar_auto_int_out_1; // @[BaseTile.scala 212:37]
  wire  intXbar_auto_int_out_2; // @[BaseTile.scala 212:37]
  wire  intXbar_auto_int_out_3; // @[BaseTile.scala 212:37]
  wire  intXbar_auto_int_out_4; // @[BaseTile.scala 212:37]
  wire [29:0] intXbar_io_covSum; // @[BaseTile.scala 212:37]
  wire  broadcast_auto_in;
  wire  broadcast_auto_out;
  wire  buffer_clock; // @[Buffer.scala 68:28]
  wire  buffer_reset; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28]
  wire [5:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28]
  wire [31:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_bufferable; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_modifiable; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_readalloc; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_writealloc; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_privileged; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_secure; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_a_bits_user_amba_prot_fetch; // @[Buffer.scala 68:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28]
  wire [5:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28]
  wire [5:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28]
  wire [31:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_bufferable; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_modifiable; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_readalloc; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_writealloc; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_privileged; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_secure; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_a_bits_user_amba_prot_fetch; // @[Buffer.scala 68:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28]
  wire [5:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire [29:0] buffer_io_covSum; // @[Buffer.scala 68:28]
  wire  fixer_clock; // @[FIFOFixer.scala 144:27]
  wire  fixer_reset; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_in_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_in_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_in_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_in_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_in_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_in_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_in_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_in_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_a_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_a_bits_size; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_out_a_bits_source; // @[FIFOFixer.scala 144:27]
  wire [31:0] fixer_auto_out_a_bits_address; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_bufferable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_modifiable; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_readalloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_writealloc; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_privileged; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_secure; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_a_bits_user_amba_prot_fetch; // @[FIFOFixer.scala 144:27]
  wire [7:0] fixer_auto_out_a_bits_mask; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_a_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_ready; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_valid; // @[FIFOFixer.scala 144:27]
  wire [2:0] fixer_auto_out_d_bits_opcode; // @[FIFOFixer.scala 144:27]
  wire [3:0] fixer_auto_out_d_bits_size; // @[FIFOFixer.scala 144:27]
  wire [5:0] fixer_auto_out_d_bits_source; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_bits_denied; // @[FIFOFixer.scala 144:27]
  wire [63:0] fixer_auto_out_d_bits_data; // @[FIFOFixer.scala 144:27]
  wire  fixer_auto_out_d_bits_corrupt; // @[FIFOFixer.scala 144:27]
  wire [29:0] fixer_io_covSum; // @[FIFOFixer.scala 144:27]
  wire  fixer_metaReset; // @[FIFOFixer.scala 144:27]
  wire  widget_auto_in_a_ready;
  wire  widget_auto_in_a_valid;
  wire [2:0] widget_auto_in_a_bits_opcode;
  wire [3:0] widget_auto_in_a_bits_size;
  wire [5:0] widget_auto_in_a_bits_source;
  wire [31:0] widget_auto_in_a_bits_address;
  wire  widget_auto_in_a_bits_user_amba_prot_bufferable;
  wire  widget_auto_in_a_bits_user_amba_prot_modifiable;
  wire  widget_auto_in_a_bits_user_amba_prot_readalloc;
  wire  widget_auto_in_a_bits_user_amba_prot_writealloc;
  wire  widget_auto_in_a_bits_user_amba_prot_privileged;
  wire  widget_auto_in_a_bits_user_amba_prot_secure;
  wire  widget_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] widget_auto_in_a_bits_mask;
  wire [63:0] widget_auto_in_a_bits_data;
  wire  widget_auto_in_d_ready;
  wire  widget_auto_in_d_valid;
  wire [2:0] widget_auto_in_d_bits_opcode;
  wire [3:0] widget_auto_in_d_bits_size;
  wire [5:0] widget_auto_in_d_bits_source;
  wire  widget_auto_in_d_bits_denied;
  wire [63:0] widget_auto_in_d_bits_data;
  wire  widget_auto_in_d_bits_corrupt;
  wire  widget_auto_out_a_ready;
  wire  widget_auto_out_a_valid;
  wire [2:0] widget_auto_out_a_bits_opcode;
  wire [3:0] widget_auto_out_a_bits_size;
  wire [5:0] widget_auto_out_a_bits_source;
  wire [31:0] widget_auto_out_a_bits_address;
  wire  widget_auto_out_a_bits_user_amba_prot_bufferable;
  wire  widget_auto_out_a_bits_user_amba_prot_modifiable;
  wire  widget_auto_out_a_bits_user_amba_prot_readalloc;
  wire  widget_auto_out_a_bits_user_amba_prot_writealloc;
  wire  widget_auto_out_a_bits_user_amba_prot_privileged;
  wire  widget_auto_out_a_bits_user_amba_prot_secure;
  wire  widget_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] widget_auto_out_a_bits_mask;
  wire [63:0] widget_auto_out_a_bits_data;
  wire  widget_auto_out_d_ready;
  wire  widget_auto_out_d_valid;
  wire [2:0] widget_auto_out_d_bits_opcode;
  wire [3:0] widget_auto_out_d_bits_size;
  wire [5:0] widget_auto_out_d_bits_source;
  wire  widget_auto_out_d_bits_denied;
  wire [63:0] widget_auto_out_d_bits_data;
  wire  widget_auto_out_d_bits_corrupt;
  wire  axi42tl_clock; // @[ToTL.scala 216:29]
  wire  axi42tl_reset; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_aw_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_aw_valid; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_in_aw_bits_id; // @[ToTL.scala 216:29]
  wire [31:0] axi42tl_auto_in_aw_bits_addr; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_in_aw_bits_len; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_aw_bits_size; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_in_aw_bits_cache; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_aw_bits_prot; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_w_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_w_valid; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_in_w_bits_data; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_in_w_bits_strb; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_w_bits_last; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_b_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_b_valid; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_in_b_bits_id; // @[ToTL.scala 216:29]
  wire [1:0] axi42tl_auto_in_b_bits_resp; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_ar_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_ar_valid; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_in_ar_bits_id; // @[ToTL.scala 216:29]
  wire [31:0] axi42tl_auto_in_ar_bits_addr; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_in_ar_bits_len; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_ar_bits_size; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_in_ar_bits_cache; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_in_ar_bits_prot; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_r_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_r_valid; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_in_r_bits_id; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_in_r_bits_data; // @[ToTL.scala 216:29]
  wire [1:0] axi42tl_auto_in_r_bits_resp; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_in_r_bits_last; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_valid; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_out_a_bits_opcode; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_out_a_bits_size; // @[ToTL.scala 216:29]
  wire [5:0] axi42tl_auto_out_a_bits_source; // @[ToTL.scala 216:29]
  wire [31:0] axi42tl_auto_out_a_bits_address; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_bufferable; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_modifiable; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_readalloc; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_writealloc; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_privileged; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_secure; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_a_bits_user_amba_prot_fetch; // @[ToTL.scala 216:29]
  wire [7:0] axi42tl_auto_out_a_bits_mask; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_out_a_bits_data; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_ready; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_valid; // @[ToTL.scala 216:29]
  wire [2:0] axi42tl_auto_out_d_bits_opcode; // @[ToTL.scala 216:29]
  wire [3:0] axi42tl_auto_out_d_bits_size; // @[ToTL.scala 216:29]
  wire [5:0] axi42tl_auto_out_d_bits_source; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_bits_denied; // @[ToTL.scala 216:29]
  wire [63:0] axi42tl_auto_out_d_bits_data; // @[ToTL.scala 216:29]
  wire  axi42tl_auto_out_d_bits_corrupt; // @[ToTL.scala 216:29]
  wire [29:0] axi42tl_io_covSum; // @[ToTL.scala 216:29]
  wire  axi42tl_metaReset; // @[ToTL.scala 216:29]
  wire  axi4yank_clock; // @[UserYanker.scala 105:30]
  wire  axi4yank_reset; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_aw_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_in_aw_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_aw_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_aw_bits_size; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_aw_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_aw_bits_prot; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_aw_bits_echo_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_w_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_w_valid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_in_w_bits_data; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_w_bits_strb; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_w_bits_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_b_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_b_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_b_bits_id; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_b_bits_resp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_b_bits_echo_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_ar_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_in_ar_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_in_ar_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_ar_bits_size; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_ar_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_in_ar_bits_prot; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_ar_bits_echo_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_in_r_bits_id; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_in_r_bits_data; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_in_r_bits_resp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_bits_echo_real_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_in_r_bits_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_aw_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_aw_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_aw_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_out_aw_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_aw_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_aw_bits_size; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_aw_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_aw_bits_prot; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_w_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_w_valid; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_out_w_bits_data; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_w_bits_strb; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_w_bits_last; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_b_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_b_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_b_bits_id; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_b_bits_resp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_ar_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_ar_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_ar_bits_id; // @[UserYanker.scala 105:30]
  wire [31:0] axi4yank_auto_out_ar_bits_addr; // @[UserYanker.scala 105:30]
  wire [7:0] axi4yank_auto_out_ar_bits_len; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_ar_bits_size; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_ar_bits_cache; // @[UserYanker.scala 105:30]
  wire [2:0] axi4yank_auto_out_ar_bits_prot; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_ready; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_valid; // @[UserYanker.scala 105:30]
  wire [3:0] axi4yank_auto_out_r_bits_id; // @[UserYanker.scala 105:30]
  wire [63:0] axi4yank_auto_out_r_bits_data; // @[UserYanker.scala 105:30]
  wire [1:0] axi4yank_auto_out_r_bits_resp; // @[UserYanker.scala 105:30]
  wire  axi4yank_auto_out_r_bits_last; // @[UserYanker.scala 105:30]
  wire [29:0] axi4yank_io_covSum; // @[UserYanker.scala 105:30]
  wire  axi4frag_clock; // @[Fragmenter.scala 205:30]
  wire  axi4frag_reset; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_aw_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_aw_valid; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_in_aw_bits_id; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_in_aw_bits_addr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_in_aw_bits_len; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_aw_bits_size; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_aw_bits_burst; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_in_aw_bits_cache; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_aw_bits_prot; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_w_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_w_valid; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_in_w_bits_data; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_in_w_bits_strb; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_w_bits_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_b_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_b_valid; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_in_b_bits_id; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_b_bits_resp; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_ar_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_ar_valid; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_in_ar_bits_id; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_in_ar_bits_addr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_in_ar_bits_len; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_ar_bits_size; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_ar_bits_burst; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_in_ar_bits_cache; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_in_ar_bits_prot; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_r_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_r_valid; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_in_r_bits_id; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_in_r_bits_data; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_in_r_bits_resp; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_in_r_bits_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_aw_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_aw_valid; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_out_aw_bits_id; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_out_aw_bits_addr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_out_aw_bits_len; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_aw_bits_size; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_out_aw_bits_cache; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_aw_bits_prot; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_aw_bits_echo_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_w_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_w_valid; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_out_w_bits_data; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_out_w_bits_strb; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_w_bits_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_b_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_b_valid; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_out_b_bits_id; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_out_b_bits_resp; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_b_bits_echo_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_ar_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_ar_valid; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_out_ar_bits_id; // @[Fragmenter.scala 205:30]
  wire [31:0] axi4frag_auto_out_ar_bits_addr; // @[Fragmenter.scala 205:30]
  wire [7:0] axi4frag_auto_out_ar_bits_len; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_ar_bits_size; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_out_ar_bits_cache; // @[Fragmenter.scala 205:30]
  wire [2:0] axi4frag_auto_out_ar_bits_prot; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_ar_bits_echo_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_r_ready; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_r_valid; // @[Fragmenter.scala 205:30]
  wire [3:0] axi4frag_auto_out_r_bits_id; // @[Fragmenter.scala 205:30]
  wire [63:0] axi4frag_auto_out_r_bits_data; // @[Fragmenter.scala 205:30]
  wire [1:0] axi4frag_auto_out_r_bits_resp; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_r_bits_echo_real_last; // @[Fragmenter.scala 205:30]
  wire  axi4frag_auto_out_r_bits_last; // @[Fragmenter.scala 205:30]
  wire [29:0] axi4frag_io_covSum; // @[Fragmenter.scala 205:30]
  wire  axi4frag_metaReset; // @[Fragmenter.scala 205:30]
  wire  core_clk_i; // @[CVA6Tile.scala 234:20]
  wire  core_rst_ni; // @[CVA6Tile.scala 234:20]
  wire [63:0] core_boot_addr_i; // @[CVA6Tile.scala 234:20]
  wire [63:0] core_hart_id_i; // @[CVA6Tile.scala 234:20]
  wire [1:0] core_irq_i; // @[CVA6Tile.scala 234:20]
  wire  core_ipi_i; // @[CVA6Tile.scala 234:20]
  wire  core_time_irq_i; // @[CVA6Tile.scala 234:20]
  wire  core_debug_req_i; // @[CVA6Tile.scala 234:20]
  wire [367:0] core_trace_o; // @[CVA6Tile.scala 234:20]
  wire  core_axi_resp_i_aw_ready; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_aw_valid; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_req_o_aw_bits_id; // @[CVA6Tile.scala 234:20]
  wire [63:0] core_axi_req_o_aw_bits_addr; // @[CVA6Tile.scala 234:20]
  wire [7:0] core_axi_req_o_aw_bits_len; // @[CVA6Tile.scala 234:20]
  wire [2:0] core_axi_req_o_aw_bits_size; // @[CVA6Tile.scala 234:20]
  wire [1:0] core_axi_req_o_aw_bits_burst; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_aw_bits_lock; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_req_o_aw_bits_cache; // @[CVA6Tile.scala 234:20]
  wire [2:0] core_axi_req_o_aw_bits_prot; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_req_o_aw_bits_qos; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_req_o_aw_bits_region; // @[CVA6Tile.scala 234:20]
  wire [5:0] core_axi_req_o_aw_bits_atop; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_aw_bits_user; // @[CVA6Tile.scala 234:20]
  wire  core_axi_resp_i_w_ready; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_w_valid; // @[CVA6Tile.scala 234:20]
  wire [63:0] core_axi_req_o_w_bits_data; // @[CVA6Tile.scala 234:20]
  wire [7:0] core_axi_req_o_w_bits_strb; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_w_bits_last; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_w_bits_user; // @[CVA6Tile.scala 234:20]
  wire  core_axi_resp_i_ar_ready; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_ar_valid; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_req_o_ar_bits_id; // @[CVA6Tile.scala 234:20]
  wire [63:0] core_axi_req_o_ar_bits_addr; // @[CVA6Tile.scala 234:20]
  wire [7:0] core_axi_req_o_ar_bits_len; // @[CVA6Tile.scala 234:20]
  wire [2:0] core_axi_req_o_ar_bits_size; // @[CVA6Tile.scala 234:20]
  wire [1:0] core_axi_req_o_ar_bits_burst; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_ar_bits_lock; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_req_o_ar_bits_cache; // @[CVA6Tile.scala 234:20]
  wire [2:0] core_axi_req_o_ar_bits_prot; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_req_o_ar_bits_qos; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_req_o_ar_bits_region; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_ar_bits_user; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_b_ready; // @[CVA6Tile.scala 234:20]
  wire  core_axi_resp_i_b_valid; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_resp_i_b_bits_id; // @[CVA6Tile.scala 234:20]
  wire [1:0] core_axi_resp_i_b_bits_resp; // @[CVA6Tile.scala 234:20]
  wire  core_axi_resp_i_b_bits_user; // @[CVA6Tile.scala 234:20]
  wire  core_axi_req_o_r_ready; // @[CVA6Tile.scala 234:20]
  wire  core_axi_resp_i_r_valid; // @[CVA6Tile.scala 234:20]
  wire [3:0] core_axi_resp_i_r_bits_id; // @[CVA6Tile.scala 234:20]
  wire [63:0] core_axi_resp_i_r_bits_data; // @[CVA6Tile.scala 234:20]
  wire [1:0] core_axi_resp_i_r_bits_resp; // @[CVA6Tile.scala 234:20]
  wire  core_axi_resp_i_r_bits_last; // @[CVA6Tile.scala 234:20]
  wire  core_axi_resp_i_r_bits_user; // @[CVA6Tile.scala 234:20]
  wire  _core_io_rst_ni_T_1 = ~reset; // @[CVA6Tile.scala 259:21]
  wire  bundleIn_0_9_4 = intXbar_auto_int_out_4; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  wire  bundleIn_0_9_3 = intXbar_auto_int_out_3; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  wire [29:0] CVA6Tile_covSum;
  wire [29:0] axi4yank_sum;
  wire [29:0] intXbar_sum;
  wire [29:0] buffer_sum;
  wire [29:0] axi4frag_sum;
  wire [29:0] fixer_sum;
  wire [29:0] axi42tl_sum;
  IntXbar_1 intXbar ( // @[BaseTile.scala 212:37]
    .auto_int_in_3_0(intXbar_auto_int_in_3_0),
    .auto_int_in_2_0(intXbar_auto_int_in_2_0),
    .auto_int_in_1_0(intXbar_auto_int_in_1_0),
    .auto_int_in_1_1(intXbar_auto_int_in_1_1),
    .auto_int_out_1(intXbar_auto_int_out_1),
    .auto_int_out_2(intXbar_auto_int_out_2),
    .auto_int_out_3(intXbar_auto_int_out_3),
    .auto_int_out_4(intXbar_auto_int_out_4),
    .io_covSum(intXbar_io_covSum)
  );
  TLBuffer_8 buffer ( // @[Buffer.scala 68:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(buffer_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(buffer_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(buffer_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(buffer_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(buffer_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(buffer_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(buffer_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(buffer_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(buffer_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(buffer_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(buffer_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(buffer_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(buffer_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(buffer_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt),
    .io_covSum(buffer_io_covSum)
  );
  TLFIFOFixer_5 fixer ( // @[FIFOFixer.scala 144:27]
    .clock(fixer_clock),
    .reset(fixer_reset),
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(fixer_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(fixer_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(fixer_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(fixer_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(fixer_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(fixer_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(fixer_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_auto_in_a_bits_data),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(fixer_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(fixer_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(fixer_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(fixer_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(fixer_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(fixer_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(fixer_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_auto_out_a_bits_data),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt),
    .io_covSum(fixer_io_covSum),
    .metaReset(fixer_metaReset)
  );
  AXI4ToTL_1 axi42tl ( // @[ToTL.scala 216:29]
    .clock(axi42tl_clock),
    .reset(axi42tl_reset),
    .auto_in_aw_ready(axi42tl_auto_in_aw_ready),
    .auto_in_aw_valid(axi42tl_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi42tl_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi42tl_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi42tl_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi42tl_auto_in_aw_bits_size),
    .auto_in_aw_bits_cache(axi42tl_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi42tl_auto_in_aw_bits_prot),
    .auto_in_w_ready(axi42tl_auto_in_w_ready),
    .auto_in_w_valid(axi42tl_auto_in_w_valid),
    .auto_in_w_bits_data(axi42tl_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi42tl_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi42tl_auto_in_w_bits_last),
    .auto_in_b_ready(axi42tl_auto_in_b_ready),
    .auto_in_b_valid(axi42tl_auto_in_b_valid),
    .auto_in_b_bits_id(axi42tl_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi42tl_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi42tl_auto_in_ar_ready),
    .auto_in_ar_valid(axi42tl_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi42tl_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi42tl_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi42tl_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi42tl_auto_in_ar_bits_size),
    .auto_in_ar_bits_cache(axi42tl_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi42tl_auto_in_ar_bits_prot),
    .auto_in_r_ready(axi42tl_auto_in_r_ready),
    .auto_in_r_valid(axi42tl_auto_in_r_valid),
    .auto_in_r_bits_id(axi42tl_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi42tl_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi42tl_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi42tl_auto_in_r_bits_last),
    .auto_out_a_ready(axi42tl_auto_out_a_ready),
    .auto_out_a_valid(axi42tl_auto_out_a_valid),
    .auto_out_a_bits_opcode(axi42tl_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(axi42tl_auto_out_a_bits_size),
    .auto_out_a_bits_source(axi42tl_auto_out_a_bits_source),
    .auto_out_a_bits_address(axi42tl_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(axi42tl_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(axi42tl_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(axi42tl_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(axi42tl_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(axi42tl_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(axi42tl_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(axi42tl_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(axi42tl_auto_out_a_bits_mask),
    .auto_out_a_bits_data(axi42tl_auto_out_a_bits_data),
    .auto_out_d_ready(axi42tl_auto_out_d_ready),
    .auto_out_d_valid(axi42tl_auto_out_d_valid),
    .auto_out_d_bits_opcode(axi42tl_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(axi42tl_auto_out_d_bits_size),
    .auto_out_d_bits_source(axi42tl_auto_out_d_bits_source),
    .auto_out_d_bits_denied(axi42tl_auto_out_d_bits_denied),
    .auto_out_d_bits_data(axi42tl_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(axi42tl_auto_out_d_bits_corrupt),
    .io_covSum(axi42tl_io_covSum),
    .metaReset(axi42tl_metaReset)
  );
  AXI4UserYanker_2 axi4yank ( // @[UserYanker.scala 105:30]
    .clock(axi4yank_clock),
    .reset(axi4yank_reset),
    .auto_in_aw_ready(axi4yank_auto_in_aw_ready),
    .auto_in_aw_valid(axi4yank_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4yank_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4yank_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4yank_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4yank_auto_in_aw_bits_size),
    .auto_in_aw_bits_cache(axi4yank_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4yank_auto_in_aw_bits_prot),
    .auto_in_aw_bits_echo_real_last(axi4yank_auto_in_aw_bits_echo_real_last),
    .auto_in_w_ready(axi4yank_auto_in_w_ready),
    .auto_in_w_valid(axi4yank_auto_in_w_valid),
    .auto_in_w_bits_data(axi4yank_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4yank_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4yank_auto_in_w_bits_last),
    .auto_in_b_ready(axi4yank_auto_in_b_ready),
    .auto_in_b_valid(axi4yank_auto_in_b_valid),
    .auto_in_b_bits_id(axi4yank_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4yank_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_real_last(axi4yank_auto_in_b_bits_echo_real_last),
    .auto_in_ar_ready(axi4yank_auto_in_ar_ready),
    .auto_in_ar_valid(axi4yank_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4yank_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4yank_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4yank_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4yank_auto_in_ar_bits_size),
    .auto_in_ar_bits_cache(axi4yank_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4yank_auto_in_ar_bits_prot),
    .auto_in_ar_bits_echo_real_last(axi4yank_auto_in_ar_bits_echo_real_last),
    .auto_in_r_ready(axi4yank_auto_in_r_ready),
    .auto_in_r_valid(axi4yank_auto_in_r_valid),
    .auto_in_r_bits_id(axi4yank_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4yank_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4yank_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_real_last(axi4yank_auto_in_r_bits_echo_real_last),
    .auto_in_r_bits_last(axi4yank_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4yank_auto_out_aw_ready),
    .auto_out_aw_valid(axi4yank_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4yank_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4yank_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4yank_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4yank_auto_out_aw_bits_size),
    .auto_out_aw_bits_cache(axi4yank_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4yank_auto_out_aw_bits_prot),
    .auto_out_w_ready(axi4yank_auto_out_w_ready),
    .auto_out_w_valid(axi4yank_auto_out_w_valid),
    .auto_out_w_bits_data(axi4yank_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4yank_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4yank_auto_out_w_bits_last),
    .auto_out_b_ready(axi4yank_auto_out_b_ready),
    .auto_out_b_valid(axi4yank_auto_out_b_valid),
    .auto_out_b_bits_id(axi4yank_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4yank_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4yank_auto_out_ar_ready),
    .auto_out_ar_valid(axi4yank_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4yank_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4yank_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4yank_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4yank_auto_out_ar_bits_size),
    .auto_out_ar_bits_cache(axi4yank_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4yank_auto_out_ar_bits_prot),
    .auto_out_r_ready(axi4yank_auto_out_r_ready),
    .auto_out_r_valid(axi4yank_auto_out_r_valid),
    .auto_out_r_bits_id(axi4yank_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4yank_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4yank_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4yank_auto_out_r_bits_last),
    .io_covSum(axi4yank_io_covSum)
  );
  AXI4Fragmenter_1 axi4frag ( // @[Fragmenter.scala 205:30]
    .clock(axi4frag_clock),
    .reset(axi4frag_reset),
    .auto_in_aw_ready(axi4frag_auto_in_aw_ready),
    .auto_in_aw_valid(axi4frag_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4frag_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4frag_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4frag_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4frag_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4frag_auto_in_aw_bits_burst),
    .auto_in_aw_bits_cache(axi4frag_auto_in_aw_bits_cache),
    .auto_in_aw_bits_prot(axi4frag_auto_in_aw_bits_prot),
    .auto_in_w_ready(axi4frag_auto_in_w_ready),
    .auto_in_w_valid(axi4frag_auto_in_w_valid),
    .auto_in_w_bits_data(axi4frag_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4frag_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4frag_auto_in_w_bits_last),
    .auto_in_b_ready(axi4frag_auto_in_b_ready),
    .auto_in_b_valid(axi4frag_auto_in_b_valid),
    .auto_in_b_bits_id(axi4frag_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4frag_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4frag_auto_in_ar_ready),
    .auto_in_ar_valid(axi4frag_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4frag_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4frag_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4frag_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4frag_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4frag_auto_in_ar_bits_burst),
    .auto_in_ar_bits_cache(axi4frag_auto_in_ar_bits_cache),
    .auto_in_ar_bits_prot(axi4frag_auto_in_ar_bits_prot),
    .auto_in_r_ready(axi4frag_auto_in_r_ready),
    .auto_in_r_valid(axi4frag_auto_in_r_valid),
    .auto_in_r_bits_id(axi4frag_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4frag_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4frag_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4frag_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4frag_auto_out_aw_ready),
    .auto_out_aw_valid(axi4frag_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4frag_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4frag_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4frag_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4frag_auto_out_aw_bits_size),
    .auto_out_aw_bits_cache(axi4frag_auto_out_aw_bits_cache),
    .auto_out_aw_bits_prot(axi4frag_auto_out_aw_bits_prot),
    .auto_out_aw_bits_echo_real_last(axi4frag_auto_out_aw_bits_echo_real_last),
    .auto_out_w_ready(axi4frag_auto_out_w_ready),
    .auto_out_w_valid(axi4frag_auto_out_w_valid),
    .auto_out_w_bits_data(axi4frag_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4frag_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4frag_auto_out_w_bits_last),
    .auto_out_b_ready(axi4frag_auto_out_b_ready),
    .auto_out_b_valid(axi4frag_auto_out_b_valid),
    .auto_out_b_bits_id(axi4frag_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4frag_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_real_last(axi4frag_auto_out_b_bits_echo_real_last),
    .auto_out_ar_ready(axi4frag_auto_out_ar_ready),
    .auto_out_ar_valid(axi4frag_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4frag_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4frag_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4frag_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4frag_auto_out_ar_bits_size),
    .auto_out_ar_bits_cache(axi4frag_auto_out_ar_bits_cache),
    .auto_out_ar_bits_prot(axi4frag_auto_out_ar_bits_prot),
    .auto_out_ar_bits_echo_real_last(axi4frag_auto_out_ar_bits_echo_real_last),
    .auto_out_r_ready(axi4frag_auto_out_r_ready),
    .auto_out_r_valid(axi4frag_auto_out_r_valid),
    .auto_out_r_bits_id(axi4frag_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4frag_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4frag_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_real_last(axi4frag_auto_out_r_bits_echo_real_last),
    .auto_out_r_bits_last(axi4frag_auto_out_r_bits_last),
    .io_covSum(axi4frag_io_covSum),
    .metaReset(axi4frag_metaReset)
  );
  CVA6CoreBlackbox
    #(.CACHE_REG_BASE_2(0), .BTB_ENTRIES(16), .CACHE_REG_SZ_2(0), .XLEN(64), .EXEC_REG_BASE_1(65536), .AXI_USER_WIDTH(1), .EXEC_REG_SZ_2(4096), .EXEC_REG_BASE_2(0), .PMP_ENTRIES(16), .EXEC_REG_SZ_0(32'd2147483648), .CACHE_REG_SZ_0(32'd2147483648), .EXEC_REG_CNT(5), .DEBUG_BASE(32'h1f800), .CACHE_REG_BASE_3(0), .EXEC_REG_SZ_1(65536), .CACHE_REG_SZ_1(0), .RAS_ENTRIES(4), .AXI_ID_WIDTH(4), .EXEC_REG_SZ_4(0), .BHT_ENTRIES(16), .EXEC_REG_BASE_3(32'h20000), .TRACEPORT_SZ(368), .CACHE_REG_BASE_4(0), .AXI_DATA_WIDTH(64), .CACHE_REG_SZ_4(0), .AXI_ADDRESS_WIDTH(64), .EXEC_REG_BASE_4(0), .CACHE_REG_BASE_1(0), .CACHE_REG_CNT(5), .CACHE_REG_SZ_3(0), .CACHE_REG_BASE_0(32'd2147483648), .EXEC_REG_BASE_0(32'd2147483648), .EXEC_REG_SZ_3(32'h2000))
    core ( // @[CVA6Tile.scala 234:20]
    .clk_i(core_clk_i),
    .rst_ni(core_rst_ni),
    .boot_addr_i(core_boot_addr_i),
    .hart_id_i(core_hart_id_i),
    .irq_i(core_irq_i),
    .ipi_i(core_ipi_i),
    .time_irq_i(core_time_irq_i),
    .debug_req_i(core_debug_req_i),
    .trace_o(core_trace_o),
    .axi_resp_i_aw_ready(core_axi_resp_i_aw_ready),
    .axi_req_o_aw_valid(core_axi_req_o_aw_valid),
    .axi_req_o_aw_bits_id(core_axi_req_o_aw_bits_id),
    .axi_req_o_aw_bits_addr(core_axi_req_o_aw_bits_addr),
    .axi_req_o_aw_bits_len(core_axi_req_o_aw_bits_len),
    .axi_req_o_aw_bits_size(core_axi_req_o_aw_bits_size),
    .axi_req_o_aw_bits_burst(core_axi_req_o_aw_bits_burst),
    .axi_req_o_aw_bits_lock(core_axi_req_o_aw_bits_lock),
    .axi_req_o_aw_bits_cache(core_axi_req_o_aw_bits_cache),
    .axi_req_o_aw_bits_prot(core_axi_req_o_aw_bits_prot),
    .axi_req_o_aw_bits_qos(core_axi_req_o_aw_bits_qos),
    .axi_req_o_aw_bits_region(core_axi_req_o_aw_bits_region),
    .axi_req_o_aw_bits_atop(core_axi_req_o_aw_bits_atop),
    .axi_req_o_aw_bits_user(core_axi_req_o_aw_bits_user),
    .axi_resp_i_w_ready(core_axi_resp_i_w_ready),
    .axi_req_o_w_valid(core_axi_req_o_w_valid),
    .axi_req_o_w_bits_data(core_axi_req_o_w_bits_data),
    .axi_req_o_w_bits_strb(core_axi_req_o_w_bits_strb),
    .axi_req_o_w_bits_last(core_axi_req_o_w_bits_last),
    .axi_req_o_w_bits_user(core_axi_req_o_w_bits_user),
    .axi_resp_i_ar_ready(core_axi_resp_i_ar_ready),
    .axi_req_o_ar_valid(core_axi_req_o_ar_valid),
    .axi_req_o_ar_bits_id(core_axi_req_o_ar_bits_id),
    .axi_req_o_ar_bits_addr(core_axi_req_o_ar_bits_addr),
    .axi_req_o_ar_bits_len(core_axi_req_o_ar_bits_len),
    .axi_req_o_ar_bits_size(core_axi_req_o_ar_bits_size),
    .axi_req_o_ar_bits_burst(core_axi_req_o_ar_bits_burst),
    .axi_req_o_ar_bits_lock(core_axi_req_o_ar_bits_lock),
    .axi_req_o_ar_bits_cache(core_axi_req_o_ar_bits_cache),
    .axi_req_o_ar_bits_prot(core_axi_req_o_ar_bits_prot),
    .axi_req_o_ar_bits_qos(core_axi_req_o_ar_bits_qos),
    .axi_req_o_ar_bits_region(core_axi_req_o_ar_bits_region),
    .axi_req_o_ar_bits_user(core_axi_req_o_ar_bits_user),
    .axi_req_o_b_ready(core_axi_req_o_b_ready),
    .axi_resp_i_b_valid(core_axi_resp_i_b_valid),
    .axi_resp_i_b_bits_id(core_axi_resp_i_b_bits_id),
    .axi_resp_i_b_bits_resp(core_axi_resp_i_b_bits_resp),
    .axi_resp_i_b_bits_user(core_axi_resp_i_b_bits_user),
    .axi_req_o_r_ready(core_axi_req_o_r_ready),
    .axi_resp_i_r_valid(core_axi_resp_i_r_valid),
    .axi_resp_i_r_bits_id(core_axi_resp_i_r_bits_id),
    .axi_resp_i_r_bits_data(core_axi_resp_i_r_bits_data),
    .axi_resp_i_r_bits_resp(core_axi_resp_i_r_bits_resp),
    .axi_resp_i_r_bits_last(core_axi_resp_i_r_bits_last),
    .axi_resp_i_r_bits_user(core_axi_resp_i_r_bits_user)
  );
  assign tlMasterXbar_auto_in_a_ready = tlMasterXbar_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_in_d_valid = tlMasterXbar_auto_out_d_valid; // @[ReadyValidCancel.scala 21:38]
  assign tlMasterXbar_auto_in_d_bits_opcode = tlMasterXbar_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_in_d_bits_size = tlMasterXbar_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_in_d_bits_source = tlMasterXbar_auto_out_d_bits_source; // @[Xbar.scala 228:69]
  assign tlMasterXbar_auto_in_d_bits_denied = tlMasterXbar_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_in_d_bits_data = tlMasterXbar_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_in_d_bits_corrupt = tlMasterXbar_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_a_valid = tlMasterXbar_auto_in_a_valid; // @[ReadyValidCancel.scala 21:38]
  assign tlMasterXbar_auto_out_a_bits_opcode = tlMasterXbar_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_param = tlMasterXbar_auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_size = tlMasterXbar_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_source = tlMasterXbar_auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign tlMasterXbar_auto_out_a_bits_address = tlMasterXbar_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_user_amba_prot_bufferable = tlMasterXbar_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_user_amba_prot_modifiable = tlMasterXbar_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_user_amba_prot_readalloc = tlMasterXbar_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_user_amba_prot_writealloc = tlMasterXbar_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_user_amba_prot_privileged = tlMasterXbar_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_user_amba_prot_secure = tlMasterXbar_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_user_amba_prot_fetch = tlMasterXbar_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_mask = tlMasterXbar_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_a_bits_data = tlMasterXbar_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tlMasterXbar_auto_out_d_ready = tlMasterXbar_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_auto_out = broadcast_auto_in; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_in_a_ready = widget_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_valid = widget_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_opcode = widget_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_size = widget_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_source = widget_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_denied = widget_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_data = widget_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_in_d_bits_corrupt = widget_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign widget_auto_out_a_valid = widget_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_opcode = widget_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_size = widget_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_source = widget_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_address = widget_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_bufferable = widget_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_modifiable = widget_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_readalloc = widget_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_writealloc = widget_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_privileged = widget_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_secure = widget_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_user_amba_prot_fetch = widget_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_mask = widget_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_a_bits_data = widget_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign widget_auto_out_d_ready = widget_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_tl_other_masters_out_a_valid = tlMasterXbar_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_opcode = tlMasterXbar_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_param = tlMasterXbar_auto_out_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_size = tlMasterXbar_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_source = tlMasterXbar_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_address = tlMasterXbar_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_user_amba_prot_bufferable =
    tlMasterXbar_auto_out_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_user_amba_prot_modifiable =
    tlMasterXbar_auto_out_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_user_amba_prot_readalloc =
    tlMasterXbar_auto_out_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_user_amba_prot_writealloc =
    tlMasterXbar_auto_out_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_user_amba_prot_privileged =
    tlMasterXbar_auto_out_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_user_amba_prot_secure = tlMasterXbar_auto_out_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_user_amba_prot_fetch = tlMasterXbar_auto_out_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_mask = tlMasterXbar_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_data = tlMasterXbar_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_d_ready = tlMasterXbar_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_valid = buffer_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_param = buffer_auto_out_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_user_amba_prot_bufferable = buffer_auto_out_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_user_amba_prot_modifiable = buffer_auto_out_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_user_amba_prot_readalloc = buffer_auto_out_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_user_amba_prot_writealloc = buffer_auto_out_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_user_amba_prot_privileged = buffer_auto_out_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_user_amba_prot_secure = buffer_auto_out_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_user_amba_prot_fetch = buffer_auto_out_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_d_ready = buffer_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_a_ready = auto_tl_other_masters_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_valid = auto_tl_other_masters_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_opcode = auto_tl_other_masters_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_size = auto_tl_other_masters_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_source = auto_tl_other_masters_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_denied = auto_tl_other_masters_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_data = auto_tl_other_masters_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_corrupt = auto_tl_other_masters_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign intXbar_auto_int_in_3_0 = auto_int_local_in_3_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intXbar_auto_int_in_2_0 = auto_int_local_in_2_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intXbar_auto_int_in_1_0 = auto_int_local_in_1_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intXbar_auto_int_in_1_1 = auto_int_local_in_1_1; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_auto_in = auto_hartid_in; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_a_valid = fixer_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_param = 3'h0; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_size = fixer_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_source = fixer_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_address = fixer_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_bufferable = fixer_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_modifiable = fixer_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_readalloc = fixer_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_writealloc = fixer_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_privileged = fixer_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_secure = fixer_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_user_amba_prot_fetch = fixer_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_a_bits_data = fixer_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign buffer_auto_in_d_ready = fixer_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign buffer_auto_out_a_ready = tlMasterXbar_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign buffer_auto_out_d_valid = tlMasterXbar_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_opcode = tlMasterXbar_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_size = tlMasterXbar_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_source = tlMasterXbar_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_denied = tlMasterXbar_auto_in_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_data = tlMasterXbar_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_corrupt = tlMasterXbar_auto_in_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign fixer_clock = clock;
  assign fixer_reset = reset;
  assign fixer_auto_in_a_valid = widget_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_size = widget_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_source = widget_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_address = widget_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_bufferable = widget_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_modifiable = widget_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_readalloc = widget_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_writealloc = widget_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_privileged = widget_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_secure = widget_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_user_amba_prot_fetch = widget_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_mask = widget_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_a_bits_data = widget_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_in_d_ready = widget_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign fixer_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_valid = axi42tl_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_opcode = axi42tl_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_size = axi42tl_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_source = axi42tl_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_address = axi42tl_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_bufferable = axi42tl_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_modifiable = axi42tl_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_readalloc = axi42tl_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_writealloc = axi42tl_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_privileged = axi42tl_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_secure = axi42tl_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_user_amba_prot_fetch = axi42tl_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_mask = axi42tl_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign widget_auto_in_a_bits_data = axi42tl_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign widget_auto_in_d_ready = axi42tl_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign widget_auto_out_a_ready = fixer_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_valid = fixer_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_size = fixer_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_source = fixer_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_denied = fixer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_data = fixer_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign widget_auto_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign axi42tl_clock = clock;
  assign axi42tl_reset = reset;
  assign axi42tl_auto_in_aw_valid = axi4yank_auto_out_aw_valid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_id = axi4yank_auto_out_aw_bits_id; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_addr = axi4yank_auto_out_aw_bits_addr; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_len = axi4yank_auto_out_aw_bits_len; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_size = axi4yank_auto_out_aw_bits_size; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_cache = axi4yank_auto_out_aw_bits_cache; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_aw_bits_prot = axi4yank_auto_out_aw_bits_prot; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_w_valid = axi4yank_auto_out_w_valid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_w_bits_data = axi4yank_auto_out_w_bits_data; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_w_bits_strb = axi4yank_auto_out_w_bits_strb; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_w_bits_last = axi4yank_auto_out_w_bits_last; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_b_ready = axi4yank_auto_out_b_ready; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_valid = axi4yank_auto_out_ar_valid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_id = axi4yank_auto_out_ar_bits_id; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_addr = axi4yank_auto_out_ar_bits_addr; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_len = axi4yank_auto_out_ar_bits_len; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_size = axi4yank_auto_out_ar_bits_size; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_cache = axi4yank_auto_out_ar_bits_cache; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_ar_bits_prot = axi4yank_auto_out_ar_bits_prot; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_in_r_ready = axi4yank_auto_out_r_ready; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_a_ready = widget_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_valid = widget_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_opcode = widget_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_size = widget_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_source = widget_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_denied = widget_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_data = widget_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign axi42tl_auto_out_d_bits_corrupt = widget_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign axi4yank_clock = clock;
  assign axi4yank_reset = reset;
  assign axi4yank_auto_in_aw_valid = axi4frag_auto_out_aw_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_id = axi4frag_auto_out_aw_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_addr = axi4frag_auto_out_aw_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_len = axi4frag_auto_out_aw_bits_len; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_size = axi4frag_auto_out_aw_bits_size; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_cache = axi4frag_auto_out_aw_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_prot = axi4frag_auto_out_aw_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_aw_bits_echo_real_last = axi4frag_auto_out_aw_bits_echo_real_last; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_valid = axi4frag_auto_out_w_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_bits_data = axi4frag_auto_out_w_bits_data; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_bits_strb = axi4frag_auto_out_w_bits_strb; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_w_bits_last = axi4frag_auto_out_w_bits_last; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_b_ready = axi4frag_auto_out_b_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_valid = axi4frag_auto_out_ar_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_id = axi4frag_auto_out_ar_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_addr = axi4frag_auto_out_ar_bits_addr; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_len = axi4frag_auto_out_ar_bits_len; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_size = axi4frag_auto_out_ar_bits_size; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_cache = axi4frag_auto_out_ar_bits_cache; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_prot = axi4frag_auto_out_ar_bits_prot; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_ar_bits_echo_real_last = axi4frag_auto_out_ar_bits_echo_real_last; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_in_r_ready = axi4frag_auto_out_r_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_aw_ready = axi42tl_auto_in_aw_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_w_ready = axi42tl_auto_in_w_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_b_valid = axi42tl_auto_in_b_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_b_bits_id = axi42tl_auto_in_b_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_b_bits_resp = axi42tl_auto_in_b_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_ar_ready = axi42tl_auto_in_ar_ready; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_valid = axi42tl_auto_in_r_valid; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_bits_id = axi42tl_auto_in_r_bits_id; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_bits_data = axi42tl_auto_in_r_bits_data; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_bits_resp = axi42tl_auto_in_r_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4yank_auto_out_r_bits_last = axi42tl_auto_in_r_bits_last; // @[LazyModule.scala 296:16]
  assign axi4frag_clock = clock;
  assign axi4frag_reset = reset;
  assign axi4frag_auto_in_aw_valid = core_axi_req_o_aw_valid; // @[Nodes.scala 1207:84 CVA6Tile.scala 287:36]
  assign axi4frag_auto_in_aw_bits_id = core_axi_req_o_aw_bits_id; // @[Nodes.scala 1207:84 CVA6Tile.scala 288:36]
  assign axi4frag_auto_in_aw_bits_addr = core_axi_req_o_aw_bits_addr[31:0]; // @[Nodes.scala 1207:84 CVA6Tile.scala 289:36]
  assign axi4frag_auto_in_aw_bits_len = core_axi_req_o_aw_bits_len; // @[Nodes.scala 1207:84 CVA6Tile.scala 290:36]
  assign axi4frag_auto_in_aw_bits_size = core_axi_req_o_aw_bits_size; // @[Nodes.scala 1207:84 CVA6Tile.scala 291:36]
  assign axi4frag_auto_in_aw_bits_burst = core_axi_req_o_aw_bits_burst; // @[Nodes.scala 1207:84 CVA6Tile.scala 292:36]
  assign axi4frag_auto_in_aw_bits_cache = core_axi_req_o_aw_bits_cache; // @[Nodes.scala 1207:84 CVA6Tile.scala 294:36]
  assign axi4frag_auto_in_aw_bits_prot = core_axi_req_o_aw_bits_prot; // @[Nodes.scala 1207:84 CVA6Tile.scala 295:36]
  assign axi4frag_auto_in_w_valid = core_axi_req_o_w_valid; // @[Nodes.scala 1207:84 CVA6Tile.scala 303:36]
  assign axi4frag_auto_in_w_bits_data = core_axi_req_o_w_bits_data; // @[Nodes.scala 1207:84 CVA6Tile.scala 304:36]
  assign axi4frag_auto_in_w_bits_strb = core_axi_req_o_w_bits_strb; // @[Nodes.scala 1207:84 CVA6Tile.scala 305:36]
  assign axi4frag_auto_in_w_bits_last = core_axi_req_o_w_bits_last; // @[Nodes.scala 1207:84 CVA6Tile.scala 306:36]
  assign axi4frag_auto_in_b_ready = core_axi_req_o_b_ready; // @[Nodes.scala 1207:84 CVA6Tile.scala 310:36]
  assign axi4frag_auto_in_ar_valid = core_axi_req_o_ar_valid; // @[Nodes.scala 1207:84 CVA6Tile.scala 317:36]
  assign axi4frag_auto_in_ar_bits_id = core_axi_req_o_ar_bits_id; // @[Nodes.scala 1207:84 CVA6Tile.scala 318:36]
  assign axi4frag_auto_in_ar_bits_addr = core_axi_req_o_ar_bits_addr[31:0]; // @[Nodes.scala 1207:84 CVA6Tile.scala 319:36]
  assign axi4frag_auto_in_ar_bits_len = core_axi_req_o_ar_bits_len; // @[Nodes.scala 1207:84 CVA6Tile.scala 320:36]
  assign axi4frag_auto_in_ar_bits_size = core_axi_req_o_ar_bits_size; // @[Nodes.scala 1207:84 CVA6Tile.scala 321:36]
  assign axi4frag_auto_in_ar_bits_burst = core_axi_req_o_ar_bits_burst; // @[Nodes.scala 1207:84 CVA6Tile.scala 322:36]
  assign axi4frag_auto_in_ar_bits_cache = core_axi_req_o_ar_bits_cache; // @[Nodes.scala 1207:84 CVA6Tile.scala 324:36]
  assign axi4frag_auto_in_ar_bits_prot = core_axi_req_o_ar_bits_prot; // @[Nodes.scala 1207:84 CVA6Tile.scala 325:36]
  assign axi4frag_auto_in_r_ready = core_axi_req_o_r_ready; // @[Nodes.scala 1207:84 CVA6Tile.scala 331:36]
  assign axi4frag_auto_out_aw_ready = axi4yank_auto_in_aw_ready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_w_ready = axi4yank_auto_in_w_ready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_b_valid = axi4yank_auto_in_b_valid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_b_bits_id = axi4yank_auto_in_b_bits_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_b_bits_resp = axi4yank_auto_in_b_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_b_bits_echo_real_last = axi4yank_auto_in_b_bits_echo_real_last; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_ar_ready = axi4yank_auto_in_ar_ready; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_valid = axi4yank_auto_in_r_valid; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_id = axi4yank_auto_in_r_bits_id; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_data = axi4yank_auto_in_r_bits_data; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_resp = axi4yank_auto_in_r_bits_resp; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_echo_real_last = axi4yank_auto_in_r_bits_echo_real_last; // @[LazyModule.scala 296:16]
  assign axi4frag_auto_out_r_bits_last = axi4yank_auto_in_r_bits_last; // @[LazyModule.scala 296:16]
  assign core_clk_i = clock; // @[CVA6Tile.scala 258:17]
  assign core_rst_ni = ~reset; // @[CVA6Tile.scala 259:21]
  assign core_boot_addr_i = 64'h80000000; // @[CVA6Tile.scala 260:23]
  assign core_hart_id_i = {{63'd0}, broadcast_auto_out}; // @[CVA6Tile.scala 261:21]
  assign core_irq_i = {bundleIn_0_9_4,bundleIn_0_9_3}; // @[Cat.scala 31:58]
  assign core_ipi_i = intXbar_auto_int_out_1; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign core_time_irq_i = intXbar_auto_int_out_2; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign core_debug_req_i = 1'h0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign core_axi_resp_i_aw_ready = axi4frag_auto_in_aw_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_w_ready = axi4frag_auto_in_w_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_ar_ready = axi4frag_auto_in_ar_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_b_valid = axi4frag_auto_in_b_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_b_bits_id = axi4frag_auto_in_b_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_b_bits_resp = axi4frag_auto_in_b_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_b_bits_user = 1'h0; // @[CVA6Tile.scala 314:36]
  assign core_axi_resp_i_r_valid = axi4frag_auto_in_r_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_r_bits_id = axi4frag_auto_in_r_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_r_bits_data = axi4frag_auto_in_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_r_bits_resp = axi4frag_auto_in_r_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_r_bits_last = axi4frag_auto_in_r_bits_last; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign core_axi_resp_i_r_bits_user = 1'h0; // @[CVA6Tile.scala 337:36]
  assign CVA6Tile_covSum = 30'h0;
  assign axi4yank_sum = CVA6Tile_covSum + axi4yank_io_covSum;
  assign intXbar_sum = axi4yank_sum + intXbar_io_covSum;
  assign buffer_sum = intXbar_sum + buffer_io_covSum;
  assign axi4frag_sum = buffer_sum + axi4frag_io_covSum;
  assign fixer_sum = axi4frag_sum + fixer_io_covSum;
  assign axi42tl_sum = fixer_sum + axi42tl_io_covSum;
  assign io_covSum = axi42tl_sum;
  assign axi4frag_metaReset = metaReset;
  assign fixer_metaReset = metaReset;
  assign axi42tl_metaReset = metaReset;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(core_axi_req_o_aw_bits_region == 4'h0) & _core_io_rst_ni_T_1) begin
          $fatal; // @[CVA6Tile.scala 298:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_core_io_rst_ni_T_1 & ~(core_axi_req_o_aw_bits_region == 4'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at CVA6Tile.scala:298 assert(core.io.axi_req_o_aw_bits_region === 0.U)\n"); // @[CVA6Tile.scala 298:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(core_axi_req_o_aw_bits_atop == 6'h0) & _core_io_rst_ni_T_1) begin
          $fatal; // @[CVA6Tile.scala 299:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_core_io_rst_ni_T_1 & ~(core_axi_req_o_aw_bits_atop == 6'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at CVA6Tile.scala:299 assert(core.io.axi_req_o_aw_bits_atop === 0.U)\n"); // @[CVA6Tile.scala 299:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~core_axi_req_o_aw_bits_user) & _core_io_rst_ni_T_1) begin
          $fatal; // @[CVA6Tile.scala 300:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_core_io_rst_ni_T_1 & ~(~core_axi_req_o_aw_bits_user)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at CVA6Tile.scala:300 assert(core.io.axi_req_o_aw_bits_user === 0.U)\n"); // @[CVA6Tile.scala 300:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~core_axi_req_o_w_bits_user) & _core_io_rst_ni_T_1) begin
          $fatal; // @[CVA6Tile.scala 308:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_core_io_rst_ni_T_1 & ~(~core_axi_req_o_w_bits_user)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at CVA6Tile.scala:308 assert(core.io.axi_req_o_w_bits_user === 0.U)\n"); // @[CVA6Tile.scala 308:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(core_axi_req_o_ar_bits_region == 4'h0) & _core_io_rst_ni_T_1) begin
          $fatal; // @[CVA6Tile.scala 328:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_core_io_rst_ni_T_1 & ~(core_axi_req_o_ar_bits_region == 4'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at CVA6Tile.scala:328 assert(core.io.axi_req_o_ar_bits_region === 0.U)\n"); // @[CVA6Tile.scala 328:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~core_axi_req_o_ar_bits_user) & _core_io_rst_ni_T_1) begin
          $fatal; // @[CVA6Tile.scala 329:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_core_io_rst_ni_T_1 & ~(~core_axi_req_o_ar_bits_user)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at CVA6Tile.scala:329 assert(core.io.axi_req_o_ar_bits_user === 0.U)\n"); // @[CVA6Tile.scala 329:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module IntSyncSyncCrossingSink(
  input         auto_in_sync_0,
  input         auto_in_sync_1,
  output        auto_out_0,
  output        auto_out_1,
  output [29:0] io_covSum
);
  wire [29:0] IntSyncSyncCrossingSink_covSum;
  assign auto_out_0 = auto_in_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_1 = auto_in_sync_1; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign IntSyncSyncCrossingSink_covSum = 30'h0;
  assign io_covSum = IntSyncSyncCrossingSink_covSum;
endmodule
module IntSyncSyncCrossingSink_1(
  input         auto_in_sync_0,
  output        auto_out_0,
  output [29:0] io_covSum
);
  wire [29:0] IntSyncSyncCrossingSink_1_covSum;
  assign auto_out_0 = auto_in_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign IntSyncSyncCrossingSink_1_covSum = 30'h0;
  assign io_covSum = IntSyncSyncCrossingSink_1_covSum;
endmodule
module AsyncResetRegVec_w1_i0(
  input         clock,
  input         reset,
  input         io_d,
  output        io_q,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  reg_; // @[AsyncResetReg.scala 64:50]
  wire [29:0] AsyncResetRegVec_w1_i0_covSum;
  assign io_q = reg_; // @[AsyncResetReg.scala 68:8]
  assign AsyncResetRegVec_w1_i0_covSum = 30'h0;
  assign io_covSum = AsyncResetRegVec_w1_i0_covSum;
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncResetReg.scala 65:16]
      reg_ <= 1'h0; // @[AsyncResetReg.scala 66:9]
    end else begin
      reg_ <= io_d; // @[AsyncResetReg.scala 64:50]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    reg_ = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IntSyncCrossingSource_1(
  input         clock,
  input         reset,
  input         auto_in_0,
  output        auto_out_sync_0,
  output [29:0] io_covSum
);
  wire  reg__clock; // @[AsyncResetReg.scala 89:21]
  wire  reg__reset; // @[AsyncResetReg.scala 89:21]
  wire  reg__io_d; // @[AsyncResetReg.scala 89:21]
  wire  reg__io_q; // @[AsyncResetReg.scala 89:21]
  wire [29:0] reg__io_covSum; // @[AsyncResetReg.scala 89:21]
  wire [29:0] IntSyncCrossingSource_1_covSum;
  wire [29:0] reg__sum;
  AsyncResetRegVec_w1_i0 reg_ ( // @[AsyncResetReg.scala 89:21]
    .clock(reg__clock),
    .reset(reg__reset),
    .io_d(reg__io_d),
    .io_q(reg__io_q),
    .io_covSum(reg__io_covSum)
  );
  assign auto_out_sync_0 = reg__io_q; // @[Crossing.scala 41:52]
  assign reg__clock = clock;
  assign reg__reset = reset;
  assign reg__io_d = auto_in_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign IntSyncCrossingSource_1_covSum = 30'h0;
  assign reg__sum = IntSyncCrossingSource_1_covSum + reg__io_covSum;
  assign io_covSum = reg__sum;
endmodule
module TilePRCIDomain(
  input         auto_tile_reset_domain_cva6_tile_hartid_in,
  output        auto_int_out_clock_xing_out_2_sync_0,
  output        auto_int_out_clock_xing_out_1_sync_0,
  output        auto_int_out_clock_xing_out_0_sync_0,
  input         auto_int_in_clock_xing_in_2_sync_0,
  input         auto_int_in_clock_xing_in_1_sync_0,
  input         auto_int_in_clock_xing_in_0_sync_0,
  input         auto_int_in_clock_xing_in_0_sync_1,
  input         auto_tl_master_clock_xing_out_a_ready,
  output        auto_tl_master_clock_xing_out_a_valid,
  output [2:0]  auto_tl_master_clock_xing_out_a_bits_opcode,
  output [2:0]  auto_tl_master_clock_xing_out_a_bits_param,
  output [3:0]  auto_tl_master_clock_xing_out_a_bits_size,
  output [5:0]  auto_tl_master_clock_xing_out_a_bits_source,
  output [31:0] auto_tl_master_clock_xing_out_a_bits_address,
  output        auto_tl_master_clock_xing_out_a_bits_user_amba_prot_bufferable,
  output        auto_tl_master_clock_xing_out_a_bits_user_amba_prot_modifiable,
  output        auto_tl_master_clock_xing_out_a_bits_user_amba_prot_readalloc,
  output        auto_tl_master_clock_xing_out_a_bits_user_amba_prot_writealloc,
  output        auto_tl_master_clock_xing_out_a_bits_user_amba_prot_privileged,
  output        auto_tl_master_clock_xing_out_a_bits_user_amba_prot_secure,
  output        auto_tl_master_clock_xing_out_a_bits_user_amba_prot_fetch,
  output [7:0]  auto_tl_master_clock_xing_out_a_bits_mask,
  output [63:0] auto_tl_master_clock_xing_out_a_bits_data,
  output        auto_tl_master_clock_xing_out_d_ready,
  input         auto_tl_master_clock_xing_out_d_valid,
  input  [2:0]  auto_tl_master_clock_xing_out_d_bits_opcode,
  input  [3:0]  auto_tl_master_clock_xing_out_d_bits_size,
  input  [5:0]  auto_tl_master_clock_xing_out_d_bits_source,
  input         auto_tl_master_clock_xing_out_d_bits_denied,
  input  [63:0] auto_tl_master_clock_xing_out_d_bits_data,
  input         auto_tl_master_clock_xing_out_d_bits_corrupt,
  input         auto_tap_clock_in_clock,
  input         auto_tap_clock_in_reset,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  tile_reset_domain_auto_cva6_tile_int_local_in_3_0;
  wire  tile_reset_domain_auto_cva6_tile_int_local_in_2_0;
  wire  tile_reset_domain_auto_cva6_tile_int_local_in_1_0;
  wire  tile_reset_domain_auto_cva6_tile_int_local_in_1_1;
  wire  tile_reset_domain_auto_cva6_tile_hartid_in;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_ready;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_valid;
  wire [2:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_opcode;
  wire [2:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_param;
  wire [3:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_size;
  wire [5:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_source;
  wire [31:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_address;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_bufferable;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_modifiable;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_readalloc;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_writealloc;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_privileged;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_secure;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_fetch;
  wire [7:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_mask;
  wire [63:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_data;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_ready;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_valid;
  wire [2:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_opcode;
  wire [3:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_size;
  wire [5:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_source;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_denied;
  wire [63:0] tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_data;
  wire  tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_corrupt;
  wire  tile_reset_domain_auto_clock_in_clock;
  wire  tile_reset_domain_auto_clock_in_reset;
  wire  tile_reset_domain_cva6_tile_clock; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_reset; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_int_local_in_3_0; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_int_local_in_2_0; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_int_local_in_1_0; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_int_local_in_1_1; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_hartid_in; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_ready; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_valid; // @[HasTiles.scala 253:53]
  wire [2:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_opcode; // @[HasTiles.scala 253:53]
  wire [2:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_param; // @[HasTiles.scala 253:53]
  wire [3:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_size; // @[HasTiles.scala 253:53]
  wire [5:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_source; // @[HasTiles.scala 253:53]
  wire [31:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_address; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_bufferable; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_modifiable; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_readalloc; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_writealloc; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_privileged; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_secure; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_fetch; // @[HasTiles.scala 253:53]
  wire [7:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_mask; // @[HasTiles.scala 253:53]
  wire [63:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_data; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_ready; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_valid; // @[HasTiles.scala 253:53]
  wire [2:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_opcode; // @[HasTiles.scala 253:53]
  wire [3:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_size; // @[HasTiles.scala 253:53]
  wire [5:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_source; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_denied; // @[HasTiles.scala 253:53]
  wire [63:0] tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_data; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_corrupt; // @[HasTiles.scala 253:53]
  wire [29:0] tile_reset_domain_cva6_tile_io_covSum; // @[HasTiles.scala 253:53]
  wire  tile_reset_domain_cva6_tile_metaReset; // @[HasTiles.scala 253:53]
  wire  clockNode_auto_in_clock;
  wire  clockNode_auto_in_reset;
  wire  clockNode_auto_out_clock;
  wire  clockNode_auto_out_reset;
  wire  buffer_auto_in_a_ready;
  wire  buffer_auto_in_a_valid;
  wire [2:0] buffer_auto_in_a_bits_opcode;
  wire [2:0] buffer_auto_in_a_bits_param;
  wire [3:0] buffer_auto_in_a_bits_size;
  wire [5:0] buffer_auto_in_a_bits_source;
  wire [31:0] buffer_auto_in_a_bits_address;
  wire  buffer_auto_in_a_bits_user_amba_prot_bufferable;
  wire  buffer_auto_in_a_bits_user_amba_prot_modifiable;
  wire  buffer_auto_in_a_bits_user_amba_prot_readalloc;
  wire  buffer_auto_in_a_bits_user_amba_prot_writealloc;
  wire  buffer_auto_in_a_bits_user_amba_prot_privileged;
  wire  buffer_auto_in_a_bits_user_amba_prot_secure;
  wire  buffer_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] buffer_auto_in_a_bits_mask;
  wire [63:0] buffer_auto_in_a_bits_data;
  wire  buffer_auto_in_d_ready;
  wire  buffer_auto_in_d_valid;
  wire [2:0] buffer_auto_in_d_bits_opcode;
  wire [3:0] buffer_auto_in_d_bits_size;
  wire [5:0] buffer_auto_in_d_bits_source;
  wire  buffer_auto_in_d_bits_denied;
  wire [63:0] buffer_auto_in_d_bits_data;
  wire  buffer_auto_in_d_bits_corrupt;
  wire  buffer_auto_out_a_ready;
  wire  buffer_auto_out_a_valid;
  wire [2:0] buffer_auto_out_a_bits_opcode;
  wire [2:0] buffer_auto_out_a_bits_param;
  wire [3:0] buffer_auto_out_a_bits_size;
  wire [5:0] buffer_auto_out_a_bits_source;
  wire [31:0] buffer_auto_out_a_bits_address;
  wire  buffer_auto_out_a_bits_user_amba_prot_bufferable;
  wire  buffer_auto_out_a_bits_user_amba_prot_modifiable;
  wire  buffer_auto_out_a_bits_user_amba_prot_readalloc;
  wire  buffer_auto_out_a_bits_user_amba_prot_writealloc;
  wire  buffer_auto_out_a_bits_user_amba_prot_privileged;
  wire  buffer_auto_out_a_bits_user_amba_prot_secure;
  wire  buffer_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] buffer_auto_out_a_bits_mask;
  wire [63:0] buffer_auto_out_a_bits_data;
  wire  buffer_auto_out_d_ready;
  wire  buffer_auto_out_d_valid;
  wire [2:0] buffer_auto_out_d_bits_opcode;
  wire [3:0] buffer_auto_out_d_bits_size;
  wire [5:0] buffer_auto_out_d_bits_source;
  wire  buffer_auto_out_d_bits_denied;
  wire [63:0] buffer_auto_out_d_bits_data;
  wire  buffer_auto_out_d_bits_corrupt;
  wire  buffer_1_clock; // @[Buffer.scala 68:28]
  wire  buffer_1_reset; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_in_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_in_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] buffer_1_auto_in_a_bits_size; // @[Buffer.scala 68:28]
  wire [5:0] buffer_1_auto_in_a_bits_source; // @[Buffer.scala 68:28]
  wire [31:0] buffer_1_auto_in_a_bits_address; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_bits_user_amba_prot_bufferable; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_bits_user_amba_prot_modifiable; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_bits_user_amba_prot_readalloc; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_bits_user_amba_prot_writealloc; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_bits_user_amba_prot_privileged; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_bits_user_amba_prot_secure; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_a_bits_user_amba_prot_fetch; // @[Buffer.scala 68:28]
  wire [7:0] buffer_1_auto_in_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_1_auto_in_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_in_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_1_auto_in_d_bits_size; // @[Buffer.scala 68:28]
  wire [5:0] buffer_1_auto_in_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_1_auto_in_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_ready; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_out_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_out_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] buffer_1_auto_out_a_bits_size; // @[Buffer.scala 68:28]
  wire [5:0] buffer_1_auto_out_a_bits_source; // @[Buffer.scala 68:28]
  wire [31:0] buffer_1_auto_out_a_bits_address; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_bits_user_amba_prot_bufferable; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_bits_user_amba_prot_modifiable; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_bits_user_amba_prot_readalloc; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_bits_user_amba_prot_writealloc; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_bits_user_amba_prot_privileged; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_bits_user_amba_prot_secure; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_a_bits_user_amba_prot_fetch; // @[Buffer.scala 68:28]
  wire [7:0] buffer_1_auto_out_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] buffer_1_auto_out_a_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_d_ready; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] buffer_1_auto_out_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] buffer_1_auto_out_d_bits_size; // @[Buffer.scala 68:28]
  wire [5:0] buffer_1_auto_out_d_bits_source; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] buffer_1_auto_out_d_bits_data; // @[Buffer.scala 68:28]
  wire  buffer_1_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire [29:0] buffer_1_io_covSum; // @[Buffer.scala 68:28]
  wire  intsink_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_auto_in_sync_1; // @[Crossing.scala 94:29]
  wire  intsink_auto_out_0; // @[Crossing.scala 94:29]
  wire  intsink_auto_out_1; // @[Crossing.scala 94:29]
  wire [29:0] intsink_io_covSum; // @[Crossing.scala 94:29]
  wire  intsink_1_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_1_auto_out_0; // @[Crossing.scala 94:29]
  wire [29:0] intsink_1_io_covSum; // @[Crossing.scala 94:29]
  wire  intsink_2_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_2_auto_out_0; // @[Crossing.scala 94:29]
  wire [29:0] intsink_2_io_covSum; // @[Crossing.scala 94:29]
  wire  intsource_1_clock; // @[Crossing.scala 26:31]
  wire  intsource_1_reset; // @[Crossing.scala 26:31]
  wire  intsource_1_auto_in_0; // @[Crossing.scala 26:31]
  wire  intsource_1_auto_out_sync_0; // @[Crossing.scala 26:31]
  wire [29:0] intsource_1_io_covSum; // @[Crossing.scala 26:31]
  wire  intsource_2_clock; // @[Crossing.scala 26:31]
  wire  intsource_2_reset; // @[Crossing.scala 26:31]
  wire  intsource_2_auto_in_0; // @[Crossing.scala 26:31]
  wire  intsource_2_auto_out_sync_0; // @[Crossing.scala 26:31]
  wire [29:0] intsource_2_io_covSum; // @[Crossing.scala 26:31]
  wire  intsource_3_clock; // @[Crossing.scala 26:31]
  wire  intsource_3_reset; // @[Crossing.scala 26:31]
  wire  intsource_3_auto_in_0; // @[Crossing.scala 26:31]
  wire  intsource_3_auto_out_sync_0; // @[Crossing.scala 26:31]
  wire [29:0] intsource_3_io_covSum; // @[Crossing.scala 26:31]
  wire [29:0] TilePRCIDomain_covSum;
  wire [29:0] tile_reset_domain_cva6_tile_sum;
  wire [29:0] intsink_2_sum;
  wire [29:0] buffer_1_sum;
  wire [29:0] intsink_sum;
  wire [29:0] intsink_1_sum;
  wire [29:0] intsource_1_sum;
  wire [29:0] intsource_2_sum;
  wire [29:0] intsource_3_sum;
  CVA6Tile tile_reset_domain_cva6_tile ( // @[HasTiles.scala 253:53]
    .clock(tile_reset_domain_cva6_tile_clock),
    .reset(tile_reset_domain_cva6_tile_reset),
    .auto_int_local_in_3_0(tile_reset_domain_cva6_tile_auto_int_local_in_3_0),
    .auto_int_local_in_2_0(tile_reset_domain_cva6_tile_auto_int_local_in_2_0),
    .auto_int_local_in_1_0(tile_reset_domain_cva6_tile_auto_int_local_in_1_0),
    .auto_int_local_in_1_1(tile_reset_domain_cva6_tile_auto_int_local_in_1_1),
    .auto_hartid_in(tile_reset_domain_cva6_tile_auto_hartid_in),
    .auto_tl_other_masters_out_a_ready(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_ready),
    .auto_tl_other_masters_out_a_valid(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_valid),
    .auto_tl_other_masters_out_a_bits_opcode(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_opcode),
    .auto_tl_other_masters_out_a_bits_param(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_param),
    .auto_tl_other_masters_out_a_bits_size(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_size),
    .auto_tl_other_masters_out_a_bits_source(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_source),
    .auto_tl_other_masters_out_a_bits_address(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_address),
    .auto_tl_other_masters_out_a_bits_user_amba_prot_bufferable(
      tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_bufferable),
    .auto_tl_other_masters_out_a_bits_user_amba_prot_modifiable(
      tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_modifiable),
    .auto_tl_other_masters_out_a_bits_user_amba_prot_readalloc(
      tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_readalloc),
    .auto_tl_other_masters_out_a_bits_user_amba_prot_writealloc(
      tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_writealloc),
    .auto_tl_other_masters_out_a_bits_user_amba_prot_privileged(
      tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_privileged),
    .auto_tl_other_masters_out_a_bits_user_amba_prot_secure(
      tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_secure),
    .auto_tl_other_masters_out_a_bits_user_amba_prot_fetch(
      tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_fetch),
    .auto_tl_other_masters_out_a_bits_mask(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_mask),
    .auto_tl_other_masters_out_a_bits_data(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_data),
    .auto_tl_other_masters_out_d_ready(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_ready),
    .auto_tl_other_masters_out_d_valid(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_valid),
    .auto_tl_other_masters_out_d_bits_opcode(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_opcode),
    .auto_tl_other_masters_out_d_bits_size(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_size),
    .auto_tl_other_masters_out_d_bits_source(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_source),
    .auto_tl_other_masters_out_d_bits_denied(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_denied),
    .auto_tl_other_masters_out_d_bits_data(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_data),
    .auto_tl_other_masters_out_d_bits_corrupt(tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_corrupt),
    .io_covSum(tile_reset_domain_cva6_tile_io_covSum),
    .metaReset(tile_reset_domain_cva6_tile_metaReset)
  );
  TLBuffer_8 buffer_1 ( // @[Buffer.scala 68:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_a_ready(buffer_1_auto_in_a_ready),
    .auto_in_a_valid(buffer_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_1_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(buffer_1_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(buffer_1_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(buffer_1_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(buffer_1_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(buffer_1_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(buffer_1_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(buffer_1_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_1_auto_in_d_ready),
    .auto_in_d_valid(buffer_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(buffer_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_1_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_1_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_1_auto_out_a_ready),
    .auto_out_a_valid(buffer_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(buffer_1_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(buffer_1_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(buffer_1_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(buffer_1_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(buffer_1_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(buffer_1_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(buffer_1_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
    .auto_out_d_ready(buffer_1_auto_out_d_ready),
    .auto_out_d_valid(buffer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
    .auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt),
    .io_covSum(buffer_1_io_covSum)
  );
  IntSyncSyncCrossingSink intsink ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_auto_in_sync_0),
    .auto_in_sync_1(intsink_auto_in_sync_1),
    .auto_out_0(intsink_auto_out_0),
    .auto_out_1(intsink_auto_out_1),
    .io_covSum(intsink_io_covSum)
  );
  IntSyncSyncCrossingSink_1 intsink_1 ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_1_auto_in_sync_0),
    .auto_out_0(intsink_1_auto_out_0),
    .io_covSum(intsink_1_io_covSum)
  );
  IntSyncSyncCrossingSink_1 intsink_2 ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_2_auto_in_sync_0),
    .auto_out_0(intsink_2_auto_out_0),
    .io_covSum(intsink_2_io_covSum)
  );
  IntSyncCrossingSource_1 intsource_1 ( // @[Crossing.scala 26:31]
    .clock(intsource_1_clock),
    .reset(intsource_1_reset),
    .auto_in_0(intsource_1_auto_in_0),
    .auto_out_sync_0(intsource_1_auto_out_sync_0),
    .io_covSum(intsource_1_io_covSum)
  );
  IntSyncCrossingSource_1 intsource_2 ( // @[Crossing.scala 26:31]
    .clock(intsource_2_clock),
    .reset(intsource_2_reset),
    .auto_in_0(intsource_2_auto_in_0),
    .auto_out_sync_0(intsource_2_auto_out_sync_0),
    .io_covSum(intsource_2_io_covSum)
  );
  IntSyncCrossingSource_1 intsource_3 ( // @[Crossing.scala 26:31]
    .clock(intsource_3_clock),
    .reset(intsource_3_reset),
    .auto_in_0(intsource_3_auto_in_0),
    .auto_out_sync_0(intsource_3_auto_out_sync_0),
    .io_covSum(intsource_3_io_covSum)
  );
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_valid =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_valid; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_opcode =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_param =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_param; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_size =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_source =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_address =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_bufferable =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_modifiable =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_readalloc =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_writealloc =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_privileged =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_secure =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_fetch =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_mask =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_data =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_ready =
    tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_ready; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_cva6_tile_clock = tile_reset_domain_auto_clock_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tile_reset_domain_cva6_tile_reset = tile_reset_domain_auto_clock_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign tile_reset_domain_cva6_tile_auto_int_local_in_3_0 = tile_reset_domain_auto_cva6_tile_int_local_in_3_0; // @[LazyModule.scala 309:16]
  assign tile_reset_domain_cva6_tile_auto_int_local_in_2_0 = tile_reset_domain_auto_cva6_tile_int_local_in_2_0; // @[LazyModule.scala 309:16]
  assign tile_reset_domain_cva6_tile_auto_int_local_in_1_0 = tile_reset_domain_auto_cva6_tile_int_local_in_1_0; // @[LazyModule.scala 309:16]
  assign tile_reset_domain_cva6_tile_auto_int_local_in_1_1 = tile_reset_domain_auto_cva6_tile_int_local_in_1_1; // @[LazyModule.scala 309:16]
  assign tile_reset_domain_cva6_tile_auto_hartid_in = tile_reset_domain_auto_cva6_tile_hartid_in; // @[LazyModule.scala 309:16]
  assign tile_reset_domain_cva6_tile_auto_tl_other_masters_out_a_ready =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_ready; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_valid =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_valid; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_opcode =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_size =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_source =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_denied =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_denied; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_data =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign tile_reset_domain_cva6_tile_auto_tl_other_masters_out_d_bits_corrupt =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign clockNode_auto_out_clock = clockNode_auto_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockNode_auto_out_reset = clockNode_auto_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_ready = buffer_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_valid = buffer_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_opcode = buffer_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_size = buffer_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_source = buffer_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_denied = buffer_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_data = buffer_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_corrupt = buffer_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_a_valid = buffer_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_opcode = buffer_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_param = buffer_auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_size = buffer_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_source = buffer_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_address = buffer_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_bufferable = buffer_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_modifiable = buffer_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_readalloc = buffer_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_writealloc = buffer_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_privileged = buffer_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_secure = buffer_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_user_amba_prot_fetch = buffer_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_mask = buffer_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_data = buffer_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_d_ready = buffer_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_int_out_clock_xing_out_2_sync_0 = intsource_3_auto_out_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_int_out_clock_xing_out_1_sync_0 = intsource_2_auto_out_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_int_out_clock_xing_out_0_sync_0 = intsource_1_auto_out_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_valid = buffer_1_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_opcode = buffer_1_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_param = buffer_1_auto_out_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_size = buffer_1_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_source = buffer_1_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_address = buffer_1_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_user_amba_prot_bufferable =
    buffer_1_auto_out_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_user_amba_prot_modifiable =
    buffer_1_auto_out_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_user_amba_prot_readalloc =
    buffer_1_auto_out_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_user_amba_prot_writealloc =
    buffer_1_auto_out_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_user_amba_prot_privileged =
    buffer_1_auto_out_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_user_amba_prot_secure = buffer_1_auto_out_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_user_amba_prot_fetch = buffer_1_auto_out_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_mask = buffer_1_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_a_bits_data = buffer_1_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_master_clock_xing_out_d_ready = buffer_1_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tile_reset_domain_auto_cva6_tile_int_local_in_3_0 = intsink_2_auto_out_0; // @[LazyModule.scala 296:16]
  assign tile_reset_domain_auto_cva6_tile_int_local_in_2_0 = intsink_1_auto_out_0; // @[LazyModule.scala 296:16]
  assign tile_reset_domain_auto_cva6_tile_int_local_in_1_0 = intsink_auto_out_0; // @[LazyModule.scala 296:16]
  assign tile_reset_domain_auto_cva6_tile_int_local_in_1_1 = intsink_auto_out_1; // @[LazyModule.scala 296:16]
  assign tile_reset_domain_auto_cva6_tile_hartid_in = auto_tile_reset_domain_cva6_tile_hartid_in; // @[LazyModule.scala 309:16]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign tile_reset_domain_auto_clock_in_clock = clockNode_auto_out_clock; // @[LazyModule.scala 296:16]
  assign tile_reset_domain_auto_clock_in_reset = clockNode_auto_out_reset; // @[LazyModule.scala 296:16]
  assign clockNode_auto_in_clock = auto_tap_clock_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign clockNode_auto_in_reset = auto_tap_clock_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_valid = tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_valid; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_opcode = tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_param = tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_param; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_size = tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_source = tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_address = tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_user_amba_prot_bufferable =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_user_amba_prot_modifiable =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_user_amba_prot_readalloc =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_user_amba_prot_writealloc =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_user_amba_prot_privileged =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_user_amba_prot_secure =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_user_amba_prot_fetch =
    tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_mask = tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_a_bits_data = tile_reset_domain_auto_cva6_tile_tl_other_masters_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign buffer_auto_in_d_ready = tile_reset_domain_auto_cva6_tile_tl_other_masters_out_d_ready; // @[LazyModule.scala 298:16]
  assign buffer_auto_out_a_ready = buffer_1_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign buffer_auto_out_d_valid = buffer_1_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_opcode = buffer_1_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_size = buffer_1_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_source = buffer_1_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_denied = buffer_1_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_data = buffer_1_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign buffer_auto_out_d_bits_corrupt = buffer_1_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign buffer_1_clock = auto_tap_clock_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_reset = auto_tap_clock_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_1_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_param = buffer_auto_out_a_bits_param; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_user_amba_prot_bufferable = buffer_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_user_amba_prot_modifiable = buffer_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_user_amba_prot_readalloc = buffer_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_user_amba_prot_writealloc = buffer_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_user_amba_prot_privileged = buffer_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_user_amba_prot_secure = buffer_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_user_amba_prot_fetch = buffer_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign buffer_1_auto_out_a_ready = auto_tl_master_clock_xing_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_out_d_valid = auto_tl_master_clock_xing_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_out_d_bits_opcode = auto_tl_master_clock_xing_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_out_d_bits_size = auto_tl_master_clock_xing_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_out_d_bits_source = auto_tl_master_clock_xing_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_out_d_bits_denied = auto_tl_master_clock_xing_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_out_d_bits_data = auto_tl_master_clock_xing_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_1_auto_out_d_bits_corrupt = auto_tl_master_clock_xing_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign intsink_auto_in_sync_0 = auto_int_in_clock_xing_in_0_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsink_auto_in_sync_1 = auto_int_in_clock_xing_in_0_sync_1; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsink_1_auto_in_sync_0 = auto_int_in_clock_xing_in_1_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsink_2_auto_in_sync_0 = auto_int_in_clock_xing_in_2_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsource_1_clock = auto_tap_clock_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsource_1_reset = auto_tap_clock_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsource_1_auto_in_0 = 1'h0; // @[LazyModule.scala 298:16]
  assign intsource_2_clock = auto_tap_clock_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsource_2_reset = auto_tap_clock_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsource_2_auto_in_0 = 1'h0; // @[LazyModule.scala 298:16]
  assign intsource_3_clock = auto_tap_clock_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsource_3_reset = auto_tap_clock_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intsource_3_auto_in_0 = 1'h0; // @[LazyModule.scala 298:16]
  assign TilePRCIDomain_covSum = 30'h0;
  assign tile_reset_domain_cva6_tile_sum = TilePRCIDomain_covSum + tile_reset_domain_cva6_tile_io_covSum;
  assign intsink_2_sum = tile_reset_domain_cva6_tile_sum + intsink_2_io_covSum;
  assign buffer_1_sum = intsink_2_sum + buffer_1_io_covSum;
  assign intsink_sum = buffer_1_sum + intsink_io_covSum;
  assign intsink_1_sum = intsink_sum + intsink_1_io_covSum;
  assign intsource_1_sum = intsink_1_sum + intsource_1_io_covSum;
  assign intsource_2_sum = intsource_1_sum + intsource_2_io_covSum;
  assign intsource_3_sum = intsource_2_sum + intsource_3_io_covSum;
  assign io_covSum = intsource_3_sum;
  assign tile_reset_domain_cva6_tile_metaReset = metaReset;
endmodule
module LevelGateway(
  input         clock,
  input         reset,
  input         io_interrupt,
  output        io_plic_valid,
  input         io_plic_ready,
  input         io_plic_complete,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  inFlight; // @[Plic.scala 34:21]
  wire  _GEN_0 = io_interrupt & io_plic_ready | inFlight; // @[Plic.scala 34:21 35:{40,51}]
  wire [29:0] LevelGateway_covSum;
  assign io_plic_valid = io_interrupt & ~inFlight; // @[Plic.scala 37:33]
  assign LevelGateway_covSum = 30'h0;
  assign io_covSum = LevelGateway_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[Plic.scala 34:21]
      inFlight <= 1'h0; // @[Plic.scala 34:21]
    end else if (io_plic_complete) begin
      inFlight <= 1'h0;
    end else begin
      inFlight <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inFlight = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PLICFanIn(
  input         io_prio_0,
  input         io_ip,
  output        io_dev,
  output        io_max,
  output [29:0] io_covSum
);
  wire [1:0] effectivePriority_1 = {io_ip,io_prio_0}; // @[Cat.scala 31:58]
  wire  _T = 2'h2 >= effectivePriority_1; // @[Plic.scala 345:20]
  wire [1:0] maxPri = _T ? 2'h2 : effectivePriority_1; // @[Misc.scala 34:9]
  wire [29:0] PLICFanIn_covSum;
  assign io_dev = _T ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  assign io_max = maxPri[0]; // @[Plic.scala 351:10]
  assign PLICFanIn_covSum = 30'h0;
  assign io_covSum = PLICFanIn_covSum;
endmodule
module Queue_33(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_read,
  input  [22:0] io_enq_bits_index,
  input  [63:0] io_enq_bits_data,
  input  [7:0]  io_enq_bits_mask,
  input  [10:0] io_enq_bits_extra_tlrr_extra_source,
  input  [1:0]  io_enq_bits_extra_tlrr_extra_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_read,
  output [22:0] io_deq_bits_index,
  output [63:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_mask,
  output [10:0] io_deq_bits_extra_tlrr_extra_source,
  output [1:0]  io_deq_bits_extra_tlrr_extra_size,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  ram_read [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_read_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_read_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_read_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_read_MPORT_en; // @[Decoupled.scala 259:95]
  reg [22:0] ram_index [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_index_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_index_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [22:0] ram_index_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [22:0] ram_index_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_index_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_index_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_index_MPORT_en; // @[Decoupled.scala 259:95]
  reg [63:0] ram_data [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 259:95]
  reg [7:0] ram_mask [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 259:95]
  reg [10:0] ram_extra_tlrr_extra_source [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_source_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [10:0] ram_extra_tlrr_extra_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [10:0] ram_extra_tlrr_extra_source_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_source_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_source_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_source_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] ram_extra_tlrr_extra_size [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_size_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [1:0] ram_extra_tlrr_extra_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_extra_tlrr_extra_size_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_size_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_size_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_extra_tlrr_extra_size_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [29:0] Queue_33_covSum;
  assign ram_read_io_deq_bits_MPORT_en = 1'h1;
  assign ram_read_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_read_io_deq_bits_MPORT_data = ram_read[ram_read_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_read_MPORT_data = io_enq_bits_read;
  assign ram_read_MPORT_addr = 1'h0;
  assign ram_read_MPORT_mask = 1'h1;
  assign ram_read_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_index_io_deq_bits_MPORT_en = 1'h1;
  assign ram_index_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_index_io_deq_bits_MPORT_data = ram_index[ram_index_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_index_MPORT_data = io_enq_bits_index;
  assign ram_index_MPORT_addr = 1'h0;
  assign ram_index_MPORT_mask = 1'h1;
  assign ram_index_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = 1'h0;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_extra_tlrr_extra_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_extra_tlrr_extra_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_extra_tlrr_extra_source_io_deq_bits_MPORT_data =
    ram_extra_tlrr_extra_source[ram_extra_tlrr_extra_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_extra_tlrr_extra_source_MPORT_data = io_enq_bits_extra_tlrr_extra_source;
  assign ram_extra_tlrr_extra_source_MPORT_addr = 1'h0;
  assign ram_extra_tlrr_extra_source_MPORT_mask = 1'h1;
  assign ram_extra_tlrr_extra_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_extra_tlrr_extra_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_extra_tlrr_extra_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_extra_tlrr_extra_size_io_deq_bits_MPORT_data =
    ram_extra_tlrr_extra_size[ram_extra_tlrr_extra_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_extra_tlrr_extra_size_MPORT_data = io_enq_bits_extra_tlrr_extra_size;
  assign ram_extra_tlrr_extra_size_MPORT_addr = 1'h0;
  assign ram_extra_tlrr_extra_size_MPORT_mask = 1'h1;
  assign ram_extra_tlrr_extra_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_read = ram_read_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_index = ram_index_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_extra_tlrr_extra_source = ram_extra_tlrr_extra_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_extra_tlrr_extra_size = ram_extra_tlrr_extra_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign Queue_33_covSum = 30'h0;
  assign io_covSum = Queue_33_covSum;
  always @(posedge clock) begin
    if (ram_read_MPORT_en & ram_read_MPORT_mask) begin
      ram_read[ram_read_MPORT_addr] <= ram_read_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_index_MPORT_en & ram_index_MPORT_mask) begin
      ram_index[ram_index_MPORT_addr] <= ram_index_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_extra_tlrr_extra_source_MPORT_en & ram_extra_tlrr_extra_source_MPORT_mask) begin
      ram_extra_tlrr_extra_source[ram_extra_tlrr_extra_source_MPORT_addr] <= ram_extra_tlrr_extra_source_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_extra_tlrr_extra_size_MPORT_en & ram_extra_tlrr_extra_size_MPORT_mask) begin
      ram_extra_tlrr_extra_size[ram_extra_tlrr_extra_size_MPORT_addr] <= ram_extra_tlrr_extra_size_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_read[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_index[initvar] = _RAND_1[22:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_extra_tlrr_extra_source[initvar] = _RAND_4[10:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_extra_tlrr_extra_size[initvar] = _RAND_5[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLPLIC(
  input         clock,
  input         reset,
  input         auto_int_in_0,
  output        auto_int_out_1_0,
  output        auto_int_out_0_0,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [1:0]  auto_in_a_bits_size,
  input  [10:0] auto_in_a_bits_source,
  input  [27:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_size,
  output [10:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  gateways_gateway_clock; // @[Plic.scala 156:27]
  wire  gateways_gateway_reset; // @[Plic.scala 156:27]
  wire  gateways_gateway_io_interrupt; // @[Plic.scala 156:27]
  wire  gateways_gateway_io_plic_valid; // @[Plic.scala 156:27]
  wire  gateways_gateway_io_plic_ready; // @[Plic.scala 156:27]
  wire  gateways_gateway_io_plic_complete; // @[Plic.scala 156:27]
  wire [29:0] gateways_gateway_io_covSum; // @[Plic.scala 156:27]
  wire  fanin_io_prio_0; // @[Plic.scala 184:25]
  wire  fanin_io_ip; // @[Plic.scala 184:25]
  wire  fanin_io_dev; // @[Plic.scala 184:25]
  wire  fanin_io_max; // @[Plic.scala 184:25]
  wire [29:0] fanin_io_covSum; // @[Plic.scala 184:25]
  wire  fanin_1_io_prio_0; // @[Plic.scala 184:25]
  wire  fanin_1_io_ip; // @[Plic.scala 184:25]
  wire  fanin_1_io_dev; // @[Plic.scala 184:25]
  wire  fanin_1_io_max; // @[Plic.scala 184:25]
  wire [29:0] fanin_1_io_covSum; // @[Plic.scala 184:25]
  wire  out_back_clock; // @[Decoupled.scala 361:21]
  wire  out_back_reset; // @[Decoupled.scala 361:21]
  wire  out_back_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  out_back_io_enq_valid; // @[Decoupled.scala 361:21]
  wire  out_back_io_enq_bits_read; // @[Decoupled.scala 361:21]
  wire [22:0] out_back_io_enq_bits_index; // @[Decoupled.scala 361:21]
  wire [63:0] out_back_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] out_back_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [10:0] out_back_io_enq_bits_extra_tlrr_extra_source; // @[Decoupled.scala 361:21]
  wire [1:0] out_back_io_enq_bits_extra_tlrr_extra_size; // @[Decoupled.scala 361:21]
  wire  out_back_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  out_back_io_deq_valid; // @[Decoupled.scala 361:21]
  wire  out_back_io_deq_bits_read; // @[Decoupled.scala 361:21]
  wire [22:0] out_back_io_deq_bits_index; // @[Decoupled.scala 361:21]
  wire [63:0] out_back_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] out_back_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [10:0] out_back_io_deq_bits_extra_tlrr_extra_source; // @[Decoupled.scala 361:21]
  wire [1:0] out_back_io_deq_bits_extra_tlrr_extra_size; // @[Decoupled.scala 361:21]
  wire [29:0] out_back_io_covSum; // @[Decoupled.scala 361:21]
  reg  priority_0; // @[Plic.scala 163:31]
  reg  threshold_0; // @[Plic.scala 166:31]
  reg  threshold_1; // @[Plic.scala 166:31]
  reg  pending_0; // @[Plic.scala 168:22]
  reg  enables_0_0; // @[Plic.scala 174:26]
  reg  enables_1_0; // @[Plic.scala 174:26]
  wire [1:0] enableVec0_0 = {enables_0_0,1'h0}; // @[Cat.scala 31:58]
  wire [1:0] enableVec0_1 = {enables_1_0,1'h0}; // @[Cat.scala 31:58]
  reg  maxDevs_0; // @[Plic.scala 181:22]
  reg  maxDevs_1; // @[Plic.scala 181:22]
  reg  bundleOut_0_0_REG; // @[Plic.scala 188:41]
  reg  bundleOut_1_0_REG; // @[Plic.scala 188:41]
  wire [3:0] out_oindex = {out_back_io_deq_bits_index[18],out_back_io_deq_bits_index[10],out_back_io_deq_bits_index[9],
    out_back_io_deq_bits_index[4]}; // @[Cat.scala 31:58]
  wire [15:0] _out_backSel_T = 16'h1 << out_oindex; // @[OneHot.scala 57:35]
  wire  out_backSel_10 = _out_backSel_T[10]; // @[RegisterRouter.scala 83:24]
  wire [22:0] out_bindex = out_back_io_deq_bits_index & 23'h7bf9ef; // @[RegisterRouter.scala 83:24]
  wire  _out_T_9 = out_bindex == 23'h0; // @[RegisterRouter.scala 83:24]
  wire  out_roready_9 = out_back_io_deq_valid & auto_in_d_ready & out_back_io_deq_bits_read & out_backSel_10 &
    out_bindex == 23'h0; // @[RegisterRouter.scala 83:24]
  wire [7:0] _out_backMask_T_23 = out_back_io_deq_bits_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_21 = out_back_io_deq_bits_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_19 = out_back_io_deq_bits_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_17 = out_back_io_deq_bits_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_15 = out_back_io_deq_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_13 = out_back_io_deq_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_11 = out_back_io_deq_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_9 = out_back_io_deq_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] out_backMask = {_out_backMask_T_23,_out_backMask_T_21,_out_backMask_T_19,_out_backMask_T_17,
    _out_backMask_T_15,_out_backMask_T_13,_out_backMask_T_11,_out_backMask_T_9}; // @[Cat.scala 31:58]
  wire  out_romask_9 = |out_backMask[63:32]; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_9 = out_roready_9 & out_romask_9; // @[RegisterRouter.scala 83:24]
  wire  out_backSel_8 = _out_backSel_T[8]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_12 = out_back_io_deq_valid & auto_in_d_ready & out_back_io_deq_bits_read & out_backSel_8 &
    out_bindex == 23'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_12 = out_roready_12 & out_romask_9; // @[RegisterRouter.scala 83:24]
  wire [1:0] _T = {out_f_roready_9,out_f_roready_12}; // @[Plic.scala 245:21]
  wire [1:0] _T_3 = _T - 2'h1; // @[Plic.scala 245:46]
  wire [1:0] _T_4 = _T & _T_3; // @[Plic.scala 245:28]
  wire  _T_7 = ~reset; // @[Plic.scala 245:11]
  wire  claiming = out_f_roready_12 & maxDevs_0 | out_f_roready_9 & maxDevs_1; // @[Plic.scala 246:96]
  wire [1:0] _claimedDevs_T = 2'h1 << claiming; // @[OneHot.scala 64:12]
  wire  claimedDevs_1 = _claimedDevs_T[1]; // @[Plic.scala 247:58]
  wire  out_woready_9 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_10 &
    out_bindex == 23'h0; // @[RegisterRouter.scala 83:24]
  wire  out_womask_9 = &out_backMask[63:32]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_9 = out_woready_9 & out_womask_9; // @[RegisterRouter.scala 83:24]
  wire  completerDev = out_back_io_deq_bits_data[32]; // @[package.scala 154:13]
  wire [1:0] _out_completer_1_T = enableVec0_1 >> completerDev; // @[Plic.scala 295:51]
  wire  completer_1 = out_f_woready_9 & _out_completer_1_T[0]; // @[Plic.scala 295:35]
  wire  out_woready_12 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_8 &
    out_bindex == 23'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_12 = out_woready_12 & out_womask_9; // @[RegisterRouter.scala 83:24]
  wire [1:0] _out_completer_0_T = enableVec0_0 >> completerDev; // @[Plic.scala 295:51]
  wire  completer_0 = out_f_woready_12 & _out_completer_0_T[0]; // @[Plic.scala 295:35]
  wire [1:0] _T_10 = {completer_1,completer_0}; // @[Plic.scala 262:23]
  wire [1:0] _T_13 = _T_10 - 2'h1; // @[Plic.scala 262:50]
  wire [1:0] _T_14 = _T_10 & _T_13; // @[Plic.scala 262:30]
  wire [1:0] _completedDevs_T_1 = 2'h1 << completerDev; // @[OneHot.scala 64:12]
  wire [1:0] completedDevs = completer_0 | completer_1 ? _completedDevs_T_1 : 2'h0; // @[Plic.scala 264:28]
  wire  out_backSel_4 = _out_backSel_T[4]; // @[RegisterRouter.scala 83:24]
  wire  out_woready_1 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_4 &
    out_bindex == 23'h0; // @[RegisterRouter.scala 83:24]
  wire  out_womask_1 = &out_backMask[1]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_1 = out_woready_1 & out_womask_1; // @[RegisterRouter.scala 83:24]
  wire  out_womask_2 = &out_backMask[32]; // @[RegisterRouter.scala 83:24]
  wire  out_backSel_0 = _out_backSel_T[0]; // @[RegisterRouter.scala 83:24]
  wire  out_woready_2 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_0 &
    out_bindex == 23'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_2 = out_woready_2 & out_womask_2; // @[RegisterRouter.scala 83:24]
  wire [32:0] out_prepend_1 = {priority_0,32'h0}; // @[Cat.scala 31:58]
  wire  out_backSel_5 = _out_backSel_T[5]; // @[RegisterRouter.scala 83:24]
  wire  out_woready_4 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_5 &
    out_bindex == 23'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_4 = out_woready_4 & out_womask_1; // @[RegisterRouter.scala 83:24]
  wire [1:0] out_prepend_3 = {pending_0,1'h0}; // @[Cat.scala 31:58]
  wire  out_womask_7 = &out_backMask[0]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_7 = out_woready_9 & out_womask_7; // @[RegisterRouter.scala 83:24]
  wire [1:0] out_prepend_4 = {1'h0,threshold_1}; // @[Cat.scala 31:58]
  wire [31:0] _out_T_99 = {{30'd0}, out_prepend_4}; // @[RegisterRouter.scala 83:24]
  wire [32:0] out_prepend_5 = {maxDevs_1,_out_T_99}; // @[Cat.scala 31:58]
  wire [63:0] _out_T_115 = {{31'd0}, out_prepend_5}; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_10 = out_woready_12 & out_womask_7; // @[RegisterRouter.scala 83:24]
  wire [1:0] out_prepend_6 = {1'h0,threshold_0}; // @[Cat.scala 31:58]
  wire [31:0] _out_T_135 = {{30'd0}, out_prepend_6}; // @[RegisterRouter.scala 83:24]
  wire [32:0] out_prepend_7 = {maxDevs_0,_out_T_135}; // @[Cat.scala 31:58]
  wire [63:0] _out_T_151 = {{31'd0}, out_prepend_7}; // @[RegisterRouter.scala 83:24]
  wire  _GEN_70 = 4'ha == out_oindex ? _out_T_9 : 1'h1; // @[MuxLiteral.scala 53:{26,32}]
  wire  _GEN_71 = 4'h8 == out_oindex ? _out_T_9 : _GEN_70; // @[MuxLiteral.scala 53:{26,32}]
  wire  _GEN_72 = 4'h5 == out_oindex ? _out_T_9 : _GEN_71; // @[MuxLiteral.scala 53:{26,32}]
  wire  _GEN_73 = 4'h4 == out_oindex ? _out_T_9 : _GEN_72; // @[MuxLiteral.scala 53:{26,32}]
  wire  _GEN_74 = 4'h2 == out_oindex ? _out_T_9 : _GEN_73; // @[MuxLiteral.scala 53:{26,32}]
  wire  out_out_bits_data_out = 4'h0 == out_oindex ? _out_T_9 : _GEN_74; // @[MuxLiteral.scala 53:{26,32}]
  wire [63:0] _GEN_76 = 4'ha == out_oindex ? _out_T_115 : 64'h0; // @[MuxLiteral.scala 53:{26,32}]
  wire [63:0] _GEN_77 = 4'h8 == out_oindex ? _out_T_151 : _GEN_76; // @[MuxLiteral.scala 53:{26,32}]
  wire [63:0] _GEN_78 = 4'h5 == out_oindex ? {{62'd0}, enableVec0_1} : _GEN_77; // @[MuxLiteral.scala 53:{26,32}]
  wire [63:0] _GEN_79 = 4'h4 == out_oindex ? {{62'd0}, enableVec0_0} : _GEN_78; // @[MuxLiteral.scala 53:{26,32}]
  wire [63:0] _GEN_80 = 4'h2 == out_oindex ? {{62'd0}, out_prepend_3} : _GEN_79; // @[MuxLiteral.scala 53:{26,32}]
  wire [63:0] out_out_bits_data_out_1 = 4'h0 == out_oindex ? {{31'd0}, out_prepend_1} : _GEN_80; // @[MuxLiteral.scala 53:{26,32}]
  wire  out_bits_read = out_back_io_deq_bits_read; // @[RegisterRouter.scala 83:{24,24}]
  reg [1:0] TLPLIC_covState; // @[Register tracking TLPLIC state]
  reg  TLPLIC_covMap [0:3]; // @[Coverage map for TLPLIC]
  wire  TLPLIC_covMap_read_en; // @[Coverage map for TLPLIC]
  wire [1:0] TLPLIC_covMap_read_addr; // @[Coverage map for TLPLIC]
  wire  TLPLIC_covMap_read_data; // @[Coverage map for TLPLIC]
  wire  TLPLIC_covMap_write_data; // @[Coverage map for TLPLIC]
  wire [1:0] TLPLIC_covMap_write_addr; // @[Coverage map for TLPLIC]
  wire  TLPLIC_covMap_write_mask; // @[Coverage map for TLPLIC]
  wire  TLPLIC_covMap_write_en; // @[Coverage map for TLPLIC]
  reg [29:0] TLPLIC_covSum; // @[Sum of coverage map]
  wire  maxDevs_0_shl;
  wire [1:0] maxDevs_0_pad;
  wire  maxDevs_1_shl;
  wire [1:0] maxDevs_1_pad;
  wire [1:0] enables_0_0_shl;
  wire [1:0] enables_0_0_pad;
  wire [1:0] enables_1_0_shl;
  wire [1:0] enables_1_0_pad;
  wire [1:0] TLPLIC_xor1;
  wire [1:0] TLPLIC_xor2;
  wire [1:0] TLPLIC_xor0;
  wire [29:0] gateways_gateway_sum;
  wire [29:0] fanin_sum;
  wire [29:0] fanin_1_sum;
  wire [29:0] out_back_sum;
  LevelGateway gateways_gateway ( // @[Plic.scala 156:27]
    .clock(gateways_gateway_clock),
    .reset(gateways_gateway_reset),
    .io_interrupt(gateways_gateway_io_interrupt),
    .io_plic_valid(gateways_gateway_io_plic_valid),
    .io_plic_ready(gateways_gateway_io_plic_ready),
    .io_plic_complete(gateways_gateway_io_plic_complete),
    .io_covSum(gateways_gateway_io_covSum)
  );
  PLICFanIn fanin ( // @[Plic.scala 184:25]
    .io_prio_0(fanin_io_prio_0),
    .io_ip(fanin_io_ip),
    .io_dev(fanin_io_dev),
    .io_max(fanin_io_max),
    .io_covSum(fanin_io_covSum)
  );
  PLICFanIn fanin_1 ( // @[Plic.scala 184:25]
    .io_prio_0(fanin_1_io_prio_0),
    .io_ip(fanin_1_io_ip),
    .io_dev(fanin_1_io_dev),
    .io_max(fanin_1_io_max),
    .io_covSum(fanin_1_io_covSum)
  );
  Queue_33 out_back ( // @[Decoupled.scala 361:21]
    .clock(out_back_clock),
    .reset(out_back_reset),
    .io_enq_ready(out_back_io_enq_ready),
    .io_enq_valid(out_back_io_enq_valid),
    .io_enq_bits_read(out_back_io_enq_bits_read),
    .io_enq_bits_index(out_back_io_enq_bits_index),
    .io_enq_bits_data(out_back_io_enq_bits_data),
    .io_enq_bits_mask(out_back_io_enq_bits_mask),
    .io_enq_bits_extra_tlrr_extra_source(out_back_io_enq_bits_extra_tlrr_extra_source),
    .io_enq_bits_extra_tlrr_extra_size(out_back_io_enq_bits_extra_tlrr_extra_size),
    .io_deq_ready(out_back_io_deq_ready),
    .io_deq_valid(out_back_io_deq_valid),
    .io_deq_bits_read(out_back_io_deq_bits_read),
    .io_deq_bits_index(out_back_io_deq_bits_index),
    .io_deq_bits_data(out_back_io_deq_bits_data),
    .io_deq_bits_mask(out_back_io_deq_bits_mask),
    .io_deq_bits_extra_tlrr_extra_source(out_back_io_deq_bits_extra_tlrr_extra_source),
    .io_deq_bits_extra_tlrr_extra_size(out_back_io_deq_bits_extra_tlrr_extra_size),
    .io_covSum(out_back_io_covSum)
  );
  assign auto_int_out_1_0 = bundleOut_1_0_REG > threshold_1; // @[Plic.scala 188:63]
  assign auto_int_out_0_0 = bundleOut_0_0_REG > threshold_0; // @[Plic.scala 188:63]
  assign auto_in_a_ready = out_back_io_enq_ready; // @[Decoupled.scala 365:17 RegisterRouter.scala 83:24]
  assign auto_in_d_valid = out_back_io_deq_valid; // @[RegisterRouter.scala 83:24]
  assign auto_in_d_bits_opcode = {{2'd0}, out_bits_read}; // @[Nodes.scala 1210:84 RegisterRouter.scala 98:19]
  assign auto_in_d_bits_size = out_back_io_deq_bits_extra_tlrr_extra_size; // @[RegisterRouter.scala 83:{24,24}]
  assign auto_in_d_bits_source = out_back_io_deq_bits_extra_tlrr_extra_source; // @[RegisterRouter.scala 83:{24,24}]
  assign auto_in_d_bits_data = out_out_bits_data_out ? out_out_bits_data_out_1 : 64'h0; // @[RegisterRouter.scala 83:24]
  assign gateways_gateway_clock = clock;
  assign gateways_gateway_reset = reset;
  assign gateways_gateway_io_interrupt = auto_int_in_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign gateways_gateway_io_plic_ready = ~pending_0; // @[Plic.scala 250:18]
  assign gateways_gateway_io_plic_complete = completedDevs[1]; // @[Plic.scala 265:33]
  assign fanin_io_prio_0 = priority_0; // @[Plic.scala 185:21]
  assign fanin_io_ip = enables_0_0 & pending_0; // @[Plic.scala 186:40]
  assign fanin_1_io_prio_0 = priority_0; // @[Plic.scala 185:21]
  assign fanin_1_io_ip = enables_1_0 & pending_0; // @[Plic.scala 186:40]
  assign out_back_clock = clock;
  assign out_back_reset = reset;
  assign out_back_io_enq_valid = auto_in_a_valid; // @[RegisterRouter.scala 83:24]
  assign out_back_io_enq_bits_read = auto_in_a_bits_opcode == 3'h4; // @[RegisterRouter.scala 72:36]
  assign out_back_io_enq_bits_index = auto_in_a_bits_address[25:3]; // @[RegisterRouter.scala 71:18 73:19]
  assign out_back_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_back_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_back_io_enq_bits_extra_tlrr_extra_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_back_io_enq_bits_extra_tlrr_extra_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_back_io_deq_ready = auto_in_d_ready; // @[RegisterRouter.scala 83:24]
  assign TLPLIC_covMap_read_en = 1'h1;
  assign TLPLIC_covMap_read_addr = TLPLIC_covState;
  assign TLPLIC_covMap_read_data = TLPLIC_covMap[TLPLIC_covMap_read_addr]; // @[Coverage map for TLPLIC]
  assign TLPLIC_covMap_write_data = 1'h1;
  assign TLPLIC_covMap_write_addr = TLPLIC_covState;
  assign TLPLIC_covMap_write_mask = 1'h1;
  assign TLPLIC_covMap_write_en = ~metaReset;
  assign maxDevs_0_shl = maxDevs_0;
  assign maxDevs_0_pad = {1'h0,maxDevs_0_shl};
  assign maxDevs_1_shl = maxDevs_1;
  assign maxDevs_1_pad = {1'h0,maxDevs_1_shl};
  assign enables_0_0_shl = {enables_0_0, 1'h0};
  assign enables_0_0_pad = enables_0_0_shl;
  assign enables_1_0_shl = {enables_1_0, 1'h0};
  assign enables_1_0_pad = enables_1_0_shl;
  assign TLPLIC_xor1 = maxDevs_0_pad ^ maxDevs_1_pad;
  assign TLPLIC_xor2 = enables_0_0_pad ^ enables_1_0_pad;
  assign TLPLIC_xor0 = TLPLIC_xor1 ^ TLPLIC_xor2;
  assign gateways_gateway_sum = TLPLIC_covSum + gateways_gateway_io_covSum;
  assign fanin_sum = gateways_gateway_sum + fanin_io_covSum;
  assign fanin_1_sum = fanin_sum + fanin_1_io_covSum;
  assign out_back_sum = fanin_1_sum + out_back_io_covSum;
  assign io_covSum = out_back_sum;
  always @(posedge clock) begin
    if (out_f_woready_2) begin // @[RegField.scala 74:88]
      priority_0 <= out_back_io_deq_bits_data[32]; // @[RegField.scala 74:92]
    end
    if (out_f_woready_10) begin // @[RegField.scala 74:88]
      threshold_0 <= out_back_io_deq_bits_data[0]; // @[RegField.scala 74:92]
    end
    if (out_f_woready_7) begin // @[RegField.scala 74:88]
      threshold_1 <= out_back_io_deq_bits_data[0]; // @[RegField.scala 74:92]
    end
    if (reset) begin // @[Plic.scala 168:22]
      pending_0 <= 1'h0; // @[Plic.scala 168:22]
    end else if (claimedDevs_1 | gateways_gateway_io_plic_valid) begin
      pending_0 <= ~claimedDevs_1;
    end
    if (out_f_woready_1) begin // @[RegField.scala 74:88]
      enables_0_0 <= out_back_io_deq_bits_data[1]; // @[RegField.scala 74:92]
    end
    if (out_f_woready_4) begin // @[RegField.scala 74:88]
      enables_1_0 <= out_back_io_deq_bits_data[1]; // @[RegField.scala 74:92]
    end
    maxDevs_0 <= fanin_io_dev; // @[Plic.scala 187:21]
    maxDevs_1 <= fanin_1_io_dev; // @[Plic.scala 187:21]
    bundleOut_0_0_REG <= fanin_io_max; // @[Plic.scala 188:41]
    bundleOut_1_0_REG <= fanin_1_io_max; // @[Plic.scala 188:41]
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_4 == 2'h0) & ~reset) begin
          $fatal; // @[Plic.scala 245:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_4 == 2'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Plic.scala:245 assert((claimer.asUInt & (claimer.asUInt - UInt(1))) === UInt(0)) // One-Hot\n"
            ); // @[Plic.scala 245:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_14 == 2'h0) & _T_7) begin
          $fatal; // @[Plic.scala 262:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & ~(_T_14 == 2'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Plic.scala:262 assert((completer.asUInt & (completer.asUInt - UInt(1))) === UInt(0)) // One-Hot\n"
            ); // @[Plic.scala 262:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(completerDev == completerDev) & _T_7) begin
          $fatal; // @[Plic.scala 292:19]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & ~(completerDev == completerDev)) begin
          $fwrite(32'h80000002,
            "Assertion failed: completerDev should be consistent for all harts\n    at Plic.scala:292 assert(completerDev === data.extract(log2Ceil(nDevices+1)-1, 0),\n"
            ); // @[Plic.scala 292:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(completerDev == completerDev) & _T_7) begin
          $fatal; // @[Plic.scala 292:19]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & ~(completerDev == completerDev)) begin
          $fwrite(32'h80000002,
            "Assertion failed: completerDev should be consistent for all harts\n    at Plic.scala:292 assert(completerDev === data.extract(log2Ceil(nDevices+1)-1, 0),\n"
            ); // @[Plic.scala 292:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    TLPLIC_covState <= TLPLIC_xor0;
    if (TLPLIC_covMap_write_en & TLPLIC_covMap_write_mask) begin
      TLPLIC_covMap[TLPLIC_covMap_write_addr] <= TLPLIC_covMap_write_data; // @[Coverage map for TLPLIC]
    end
    if (!(TLPLIC_covMap_read_data | metaReset)) begin
      TLPLIC_covSum <= TLPLIC_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    TLPLIC_covMap[initvar] = 0; //_11[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  priority_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  threshold_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  threshold_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pending_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  enables_0_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  enables_1_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  maxDevs_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  maxDevs_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  bundleOut_0_0_REG = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  bundleOut_1_0_REG = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  TLPLIC_covState = 0; //_10[1:0];
  _RAND_12 = {1{`RANDOM}};
  TLPLIC_covSum = 0; //_12[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain(
  input         auto_plic_int_in_0,
  output        auto_plic_int_out_1_0,
  output        auto_plic_int_out_0_0,
  output        auto_plic_in_a_ready,
  input         auto_plic_in_a_valid,
  input  [2:0]  auto_plic_in_a_bits_opcode,
  input  [1:0]  auto_plic_in_a_bits_size,
  input  [10:0] auto_plic_in_a_bits_source,
  input  [27:0] auto_plic_in_a_bits_address,
  input  [7:0]  auto_plic_in_a_bits_mask,
  input  [63:0] auto_plic_in_a_bits_data,
  input         auto_plic_in_d_ready,
  output        auto_plic_in_d_valid,
  output [2:0]  auto_plic_in_d_bits_opcode,
  output [1:0]  auto_plic_in_d_bits_size,
  output [10:0] auto_plic_in_d_bits_source,
  output [63:0] auto_plic_in_d_bits_data,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  plic_clock; // @[Plic.scala 362:46]
  wire  plic_reset; // @[Plic.scala 362:46]
  wire  plic_auto_int_in_0; // @[Plic.scala 362:46]
  wire  plic_auto_int_out_1_0; // @[Plic.scala 362:46]
  wire  plic_auto_int_out_0_0; // @[Plic.scala 362:46]
  wire  plic_auto_in_a_ready; // @[Plic.scala 362:46]
  wire  plic_auto_in_a_valid; // @[Plic.scala 362:46]
  wire [2:0] plic_auto_in_a_bits_opcode; // @[Plic.scala 362:46]
  wire [1:0] plic_auto_in_a_bits_size; // @[Plic.scala 362:46]
  wire [10:0] plic_auto_in_a_bits_source; // @[Plic.scala 362:46]
  wire [27:0] plic_auto_in_a_bits_address; // @[Plic.scala 362:46]
  wire [7:0] plic_auto_in_a_bits_mask; // @[Plic.scala 362:46]
  wire [63:0] plic_auto_in_a_bits_data; // @[Plic.scala 362:46]
  wire  plic_auto_in_d_ready; // @[Plic.scala 362:46]
  wire  plic_auto_in_d_valid; // @[Plic.scala 362:46]
  wire [2:0] plic_auto_in_d_bits_opcode; // @[Plic.scala 362:46]
  wire [1:0] plic_auto_in_d_bits_size; // @[Plic.scala 362:46]
  wire [10:0] plic_auto_in_d_bits_source; // @[Plic.scala 362:46]
  wire [63:0] plic_auto_in_d_bits_data; // @[Plic.scala 362:46]
  wire [29:0] plic_io_covSum; // @[Plic.scala 362:46]
  wire  plic_metaReset; // @[Plic.scala 362:46]
  wire [29:0] ClockSinkDomain_covSum;
  wire [29:0] plic_sum;
  TLPLIC plic ( // @[Plic.scala 362:46]
    .clock(plic_clock),
    .reset(plic_reset),
    .auto_int_in_0(plic_auto_int_in_0),
    .auto_int_out_1_0(plic_auto_int_out_1_0),
    .auto_int_out_0_0(plic_auto_int_out_0_0),
    .auto_in_a_ready(plic_auto_in_a_ready),
    .auto_in_a_valid(plic_auto_in_a_valid),
    .auto_in_a_bits_opcode(plic_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(plic_auto_in_a_bits_size),
    .auto_in_a_bits_source(plic_auto_in_a_bits_source),
    .auto_in_a_bits_address(plic_auto_in_a_bits_address),
    .auto_in_a_bits_mask(plic_auto_in_a_bits_mask),
    .auto_in_a_bits_data(plic_auto_in_a_bits_data),
    .auto_in_d_ready(plic_auto_in_d_ready),
    .auto_in_d_valid(plic_auto_in_d_valid),
    .auto_in_d_bits_opcode(plic_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(plic_auto_in_d_bits_size),
    .auto_in_d_bits_source(plic_auto_in_d_bits_source),
    .auto_in_d_bits_data(plic_auto_in_d_bits_data),
    .io_covSum(plic_io_covSum),
    .metaReset(plic_metaReset)
  );
  assign auto_plic_int_out_1_0 = plic_auto_int_out_1_0; // @[LazyModule.scala 311:12]
  assign auto_plic_int_out_0_0 = plic_auto_int_out_0_0; // @[LazyModule.scala 311:12]
  assign auto_plic_in_a_ready = plic_auto_in_a_ready; // @[LazyModule.scala 309:16]
  assign auto_plic_in_d_valid = plic_auto_in_d_valid; // @[LazyModule.scala 309:16]
  assign auto_plic_in_d_bits_opcode = plic_auto_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign auto_plic_in_d_bits_size = plic_auto_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_plic_in_d_bits_source = plic_auto_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign auto_plic_in_d_bits_data = plic_auto_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign plic_clock = auto_clock_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign plic_reset = auto_clock_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign plic_auto_int_in_0 = auto_plic_int_in_0; // @[LazyModule.scala 309:16]
  assign plic_auto_in_a_valid = auto_plic_in_a_valid; // @[LazyModule.scala 309:16]
  assign plic_auto_in_a_bits_opcode = auto_plic_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign plic_auto_in_a_bits_size = auto_plic_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign plic_auto_in_a_bits_source = auto_plic_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign plic_auto_in_a_bits_address = auto_plic_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign plic_auto_in_a_bits_mask = auto_plic_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign plic_auto_in_a_bits_data = auto_plic_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign plic_auto_in_d_ready = auto_plic_in_d_ready; // @[LazyModule.scala 309:16]
  assign ClockSinkDomain_covSum = 30'h0;
  assign plic_sum = ClockSinkDomain_covSum + plic_io_covSum;
  assign io_covSum = plic_sum;
  assign plic_metaReset = metaReset;
endmodule
module CLINT(
  input         clock,
  input         reset,
  output        auto_int_out_0,
  output        auto_int_out_1,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [1:0]  auto_in_a_bits_size,
  input  [10:0] auto_in_a_bits_source,
  input  [25:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_size,
  output [10:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input         io_rtcTick,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] time_; // @[CLINT.scala 69:23]
  wire [63:0] _time_T_1 = time_ + 64'h1; // @[CLINT.scala 70:38]
  reg [63:0] timecmp_0; // @[CLINT.scala 73:41]
  reg  ipi_0; // @[CLINT.scala 74:41]
  wire [7:0] oldBytes__0 = timecmp_0[7:0]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes__1 = timecmp_0[15:8]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes__2 = timecmp_0[23:16]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes__3 = timecmp_0[31:24]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes__4 = timecmp_0[39:32]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes__5 = timecmp_0[47:40]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes__6 = timecmp_0[55:48]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes__7 = timecmp_0[63:56]; // @[RegField.scala 151:53]
  wire  in_bits_read = auto_in_a_bits_opcode == 3'h4; // @[RegisterRouter.scala 72:36]
  wire [12:0] in_bits_index = auto_in_a_bits_address[15:3]; // @[RegisterRouter.scala 71:18 73:19]
  wire [1:0] out_iindex = {in_bits_index[12],in_bits_index[11]}; // @[Cat.scala 31:58]
  wire [12:0] out_findex = in_bits_index & 13'h7ff; // @[RegisterRouter.scala 83:24]
  wire  _out_T_4 = out_findex == 13'h7ff; // @[RegisterRouter.scala 83:24]
  wire  _out_T_2 = out_findex == 13'h0; // @[RegisterRouter.scala 83:24]
  wire [3:0] _out_backSel_T = 4'h1 << out_iindex; // @[OneHot.scala 57:35]
  wire  out_backSel_1 = _out_backSel_T[1]; // @[RegisterRouter.scala 83:24]
  wire  out_woready_2 = auto_in_a_valid & auto_in_d_ready & ~in_bits_read & out_backSel_1 & out_findex == 13'h0; // @[RegisterRouter.scala 83:24]
  wire [7:0] _out_backMask_T_23 = auto_in_a_bits_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_21 = auto_in_a_bits_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_19 = auto_in_a_bits_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_17 = auto_in_a_bits_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_15 = auto_in_a_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_13 = auto_in_a_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_11 = auto_in_a_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_9 = auto_in_a_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] out_backMask = {_out_backMask_T_23,_out_backMask_T_21,_out_backMask_T_19,_out_backMask_T_17,
    _out_backMask_T_15,_out_backMask_T_13,_out_backMask_T_11,_out_backMask_T_9}; // @[Cat.scala 31:58]
  wire  out_womask_2 = &out_backMask[7:0]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_2 = out_woready_2 & out_womask_2; // @[RegisterRouter.scala 83:24]
  wire  out_womask_3 = &out_backMask[15:8]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_3 = out_woready_2 & out_womask_3; // @[RegisterRouter.scala 83:24]
  wire  out_womask_4 = &out_backMask[23:16]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_4 = out_woready_2 & out_womask_4; // @[RegisterRouter.scala 83:24]
  wire  out_womask_5 = &out_backMask[31:24]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_5 = out_woready_2 & out_womask_5; // @[RegisterRouter.scala 83:24]
  wire  out_womask_6 = &out_backMask[39:32]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_6 = out_woready_2 & out_womask_6; // @[RegisterRouter.scala 83:24]
  wire  out_womask_7 = &out_backMask[47:40]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_7 = out_woready_2 & out_womask_7; // @[RegisterRouter.scala 83:24]
  wire  out_womask_8 = &out_backMask[55:48]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_8 = out_woready_2 & out_womask_8; // @[RegisterRouter.scala 83:24]
  wire  out_womask_9 = &out_backMask[63:56]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_9 = out_woready_2 & out_womask_9; // @[RegisterRouter.scala 83:24]
  wire [7:0] newBytes__1 = out_f_woready_3 ? auto_in_a_bits_data[15:8] : oldBytes__1; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes__0 = out_f_woready_2 ? auto_in_a_bits_data[7:0] : oldBytes__0; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes__3 = out_f_woready_5 ? auto_in_a_bits_data[31:24] : oldBytes__3; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes__2 = out_f_woready_4 ? auto_in_a_bits_data[23:16] : oldBytes__2; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes__5 = out_f_woready_7 ? auto_in_a_bits_data[47:40] : oldBytes__5; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes__4 = out_f_woready_6 ? auto_in_a_bits_data[39:32] : oldBytes__4; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes__7 = out_f_woready_9 ? auto_in_a_bits_data[63:56] : oldBytes__7; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes__6 = out_f_woready_8 ? auto_in_a_bits_data[55:48] : oldBytes__6; // @[RegField.scala 158:{20,33}]
  wire [63:0] _timecmp_0_T = {newBytes__7,newBytes__6,newBytes__5,newBytes__4,newBytes__3,newBytes__2,newBytes__1,
    newBytes__0}; // @[RegField.scala 154:52]
  wire [7:0] oldBytes_1_0 = time_[7:0]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes_1_1 = time_[15:8]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes_1_2 = time_[23:16]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes_1_3 = time_[31:24]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes_1_4 = time_[39:32]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes_1_5 = time_[47:40]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes_1_6 = time_[55:48]; // @[RegField.scala 151:53]
  wire [7:0] oldBytes_1_7 = time_[63:56]; // @[RegField.scala 151:53]
  wire  out_backSel_2 = _out_backSel_T[2]; // @[RegisterRouter.scala 83:24]
  wire  out_woready_10 = auto_in_a_valid & auto_in_d_ready & ~in_bits_read & out_backSel_2 & out_findex == 13'h7ff; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_10 = out_woready_10 & out_womask_2; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_11 = out_woready_10 & out_womask_3; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_12 = out_woready_10 & out_womask_4; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_13 = out_woready_10 & out_womask_5; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_14 = out_woready_10 & out_womask_6; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_15 = out_woready_10 & out_womask_7; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_16 = out_woready_10 & out_womask_8; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_17 = out_woready_10 & out_womask_9; // @[RegisterRouter.scala 83:24]
  wire [7:0] newBytes_1_1 = out_f_woready_11 ? auto_in_a_bits_data[15:8] : oldBytes_1_1; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes_1_0 = out_f_woready_10 ? auto_in_a_bits_data[7:0] : oldBytes_1_0; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes_1_3 = out_f_woready_13 ? auto_in_a_bits_data[31:24] : oldBytes_1_3; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes_1_2 = out_f_woready_12 ? auto_in_a_bits_data[23:16] : oldBytes_1_2; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes_1_5 = out_f_woready_15 ? auto_in_a_bits_data[47:40] : oldBytes_1_5; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes_1_4 = out_f_woready_14 ? auto_in_a_bits_data[39:32] : oldBytes_1_4; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes_1_7 = out_f_woready_17 ? auto_in_a_bits_data[63:56] : oldBytes_1_7; // @[RegField.scala 158:{20,33}]
  wire [7:0] newBytes_1_6 = out_f_woready_16 ? auto_in_a_bits_data[55:48] : oldBytes_1_6; // @[RegField.scala 158:{20,33}]
  wire [63:0] _time_T_2 = {newBytes_1_7,newBytes_1_6,newBytes_1_5,newBytes_1_4,newBytes_1_3,newBytes_1_2,newBytes_1_1,
    newBytes_1_0}; // @[RegField.scala 154:52]
  wire  out_womask = &out_backMask[0]; // @[RegisterRouter.scala 83:24]
  wire  out_backSel_0 = _out_backSel_T[0]; // @[RegisterRouter.scala 83:24]
  wire  out_woready_0 = auto_in_a_valid & auto_in_d_ready & ~in_bits_read & out_backSel_0 & out_findex == 13'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready = out_woready_0 & out_womask; // @[RegisterRouter.scala 83:24]
  wire [1:0] out_prepend = {1'h0,ipi_0}; // @[Cat.scala 31:58]
  wire [31:0] _out_T_24 = {{30'd0}, out_prepend}; // @[RegisterRouter.scala 83:24]
  wire [63:0] out_prepend_7 = {oldBytes__7,oldBytes__6,oldBytes__5,oldBytes__4,oldBytes__3,oldBytes__2,oldBytes__1,
    oldBytes__0}; // @[Cat.scala 31:58]
  wire [63:0] out_prepend_14 = {oldBytes_1_7,oldBytes_1_6,oldBytes_1_5,oldBytes_1_4,oldBytes_1_3,oldBytes_1_2,
    oldBytes_1_1,oldBytes_1_0}; // @[Cat.scala 31:58]
  wire  _GEN_37 = 2'h1 == out_iindex ? _out_T_2 : _out_T_2; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_38 = 2'h2 == out_iindex ? _out_T_4 : _GEN_37; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_39 = 2'h3 == out_iindex | _GEN_38; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _out_out_bits_data_WIRE_1_0 = {{32'd0}, _out_T_24}; // @[MuxLiteral.scala 48:{48,48}]
  wire [63:0] _GEN_41 = 2'h1 == out_iindex ? out_prepend_7 : _out_out_bits_data_WIRE_1_0; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_42 = 2'h2 == out_iindex ? out_prepend_14 : _GEN_41; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_43 = 2'h3 == out_iindex ? 64'h0 : _GEN_42; // @[MuxLiteral.scala 48:{10,10}]
  wire [29:0] CLINT_covSum;
  assign auto_int_out_0 = ipi_0; // @[CLINT.scala 78:37]
  assign auto_int_out_1 = time_ >= timecmp_0; // @[CLINT.scala 79:43]
  assign auto_in_a_ready = auto_in_d_ready; // @[RegisterRouter.scala 83:24]
  assign auto_in_d_valid = auto_in_a_valid; // @[RegisterRouter.scala 83:24]
  assign auto_in_d_bits_opcode = {{2'd0}, in_bits_read}; // @[Nodes.scala 1210:84 RegisterRouter.scala 98:19]
  assign auto_in_d_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_in_d_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_in_d_bits_data = _GEN_39 ? _GEN_43 : 64'h0; // @[RegisterRouter.scala 83:24]
  assign CLINT_covSum = 30'h0;
  assign io_covSum = CLINT_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[CLINT.scala 69:23]
      time_ <= 64'h0; // @[CLINT.scala 69:23]
    end else if (out_f_woready_10 | out_f_woready_11 | out_f_woready_12 | out_f_woready_13 | out_f_woready_14 |
      out_f_woready_15 | out_f_woready_16 | out_f_woready_17) begin
      time_ <= _time_T_2;
    end else if (io_rtcTick) begin
      time_ <= _time_T_1;
    end
    if (out_f_woready_2 | out_f_woready_3 | out_f_woready_4 | out_f_woready_5 | out_f_woready_6 | out_f_woready_7 |
      out_f_woready_8 | out_f_woready_9) begin // @[RegField.scala 154:34]
      timecmp_0 <= _timecmp_0_T; // @[RegField.scala 154:40]
    end
    if (reset) begin // @[CLINT.scala 74:41]
      ipi_0 <= 1'h0; // @[CLINT.scala 74:41]
    end else if (out_f_woready) begin
      ipi_0 <= auto_in_a_bits_data[0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  time_ = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  timecmp_0 = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  ipi_0 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BundleBridgeNexus_15(
  output        auto_out,
  output [29:0] io_covSum
);
  wire  outputs_0 = 1'h0; // @[HasTiles.scala 162:32]
  wire [29:0] BundleBridgeNexus_15_covSum;
  assign auto_out = outputs_0; // @[Nodes.scala 1207:84 BundleBridge.scala 151:67]
  assign BundleBridgeNexus_15_covSum = 30'h0;
  assign io_covSum = BundleBridgeNexus_15_covSum;
endmodule
module AsyncResetRegVec_w2_i0(
  input         clock,
  input         reset,
  input  [1:0]  io_d,
  output [1:0]  io_q,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] reg_; // @[AsyncResetReg.scala 64:50]
  wire [29:0] AsyncResetRegVec_w2_i0_covSum;
  assign io_q = reg_; // @[AsyncResetReg.scala 68:8]
  assign AsyncResetRegVec_w2_i0_covSum = 30'h0;
  assign io_covSum = AsyncResetRegVec_w2_i0_covSum;
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncResetReg.scala 65:16]
      reg_ <= 2'h0; // @[AsyncResetReg.scala 66:9]
    end else begin
      reg_ <= io_d; // @[AsyncResetReg.scala 64:50]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    reg_ = 2'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IntSyncCrossingSource_4(
  input         clock,
  input         reset,
  input         auto_in_0,
  input         auto_in_1,
  output        auto_out_sync_0,
  output        auto_out_sync_1,
  output [29:0] io_covSum
);
  wire  reg__clock; // @[AsyncResetReg.scala 89:21]
  wire  reg__reset; // @[AsyncResetReg.scala 89:21]
  wire [1:0] reg__io_d; // @[AsyncResetReg.scala 89:21]
  wire [1:0] reg__io_q; // @[AsyncResetReg.scala 89:21]
  wire [29:0] reg__io_covSum; // @[AsyncResetReg.scala 89:21]
  wire [29:0] IntSyncCrossingSource_4_covSum;
  wire [29:0] reg__sum;
  AsyncResetRegVec_w2_i0 reg_ ( // @[AsyncResetReg.scala 89:21]
    .clock(reg__clock),
    .reset(reg__reset),
    .io_d(reg__io_d),
    .io_q(reg__io_q),
    .io_covSum(reg__io_covSum)
  );
  assign auto_out_sync_0 = reg__io_q[0]; // @[Crossing.scala 41:52]
  assign auto_out_sync_1 = reg__io_q[1]; // @[Crossing.scala 41:52]
  assign reg__clock = clock;
  assign reg__reset = reset;
  assign reg__io_d = {auto_in_1,auto_in_0}; // @[Cat.scala 31:58]
  assign IntSyncCrossingSource_4_covSum = 30'h0;
  assign reg__sum = IntSyncCrossingSource_4_covSum + reg__io_covSum;
  assign io_covSum = reg__sum;
endmodule
module TLROM(
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [1:0]  auto_in_a_bits_size,
  input  [10:0] auto_in_a_bits_source,
  input  [16:0] auto_in_a_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [1:0]  auto_in_d_bits_size,
  output [10:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  output [29:0] io_covSum
);
  wire [8:0] index = auto_in_a_bits_address[11:3]; // @[BootROM.scala 49:34]
  wire [3:0] high = auto_in_a_bits_address[15:12]; // @[BootROM.scala 50:68]
  wire [63:0] _GEN_1 = 9'h1 == index ? 64'h84024581f1402573 : 64'h204377c105073; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_2 = 9'h2 == index ? 64'h82090000edfe0dd0 : _GEN_1; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_3 = 9'h3 == index ? 64'h8407000038000000 : _GEN_2; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_4 = 9'h4 == index ? 64'h1100000028000000 : _GEN_3; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_5 = 9'h5 == index ? 64'h10000000 : _GEN_4; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_6 = 9'h6 == index ? 64'h4c070000fe010000 : _GEN_5; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_7 = 9'h7 == index ? 64'h0 : _GEN_6; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_8 = 9'h8 == index ? 64'h0 : _GEN_7; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_9 = 9'h9 == index ? 64'h1000000 : _GEN_8; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_10 = 9'ha == index ? 64'h400000003000000 : _GEN_9; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_11 = 9'hb == index ? 64'h100000000000000 : _GEN_10; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_12 = 9'hc == index ? 64'h400000003000000 : _GEN_11; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_13 = 9'hd == index ? 64'h10000000f000000 : _GEN_12; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_14 = 9'he == index ? 64'h1100000003000000 : _GEN_13; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_15 = 9'hf == index ? 64'h2c766a7a1b000000 : _GEN_14; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_16 = 9'h10 == index ? 64'h7069687372617473 : _GEN_15; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_17 = 9'h11 == index ? 64'h7665642d : _GEN_16; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_18 = 9'h12 == index ? 64'hd00000003000000 : _GEN_17; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_19 = 9'h13 == index ? 64'h2c766a7a26000000 : _GEN_18; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_20 = 9'h14 == index ? 64'h7069687372617473 : _GEN_19; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_21 = 9'h15 == index ? 64'h100000000000000 : _GEN_20; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_22 = 9'h16 == index ? 64'h73657361696c61 : _GEN_21; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_23 = 9'h17 == index ? 64'h1500000003000000 : _GEN_22; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_24 = 9'h18 == index ? 64'h636f732f2c000000 : _GEN_23; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_25 = 9'h19 == index ? 64'h406c61697265732f : _GEN_24; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_26 = 9'h1a == index ? 64'h3030303030303436 : _GEN_25; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_27 = 9'h1b == index ? 64'h200000000000000 : _GEN_26; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_28 = 9'h1c == index ? 64'h736f686301000000 : _GEN_27; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_29 = 9'h1d == index ? 64'h300000000006e65 : _GEN_28; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_30 = 9'h1e == index ? 64'h3400000008000000 : _GEN_29; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_31 = 9'h1f == index ? 64'h726c73616b6f6e : _GEN_30; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_32 = 9'h20 == index ? 64'h100000002000000 : _GEN_31; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_33 = 9'h21 == index ? 64'h73757063 : _GEN_32; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_34 = 9'h22 == index ? 64'h400000003000000 : _GEN_33; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_35 = 9'h23 == index ? 64'h100000000000000 : _GEN_34; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_36 = 9'h24 == index ? 64'h400000003000000 : _GEN_35; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_37 = 9'h25 == index ? 64'hf000000 : _GEN_36; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_38 = 9'h26 == index ? 64'h400000003000000 : _GEN_37; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_39 = 9'h27 == index ? 64'h40420f003d000000 : _GEN_38; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_40 = 9'h28 == index ? 64'h4075706301000000 : _GEN_39; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_41 = 9'h29 == index ? 64'h300000000000030 : _GEN_40; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_42 = 9'h2a == index ? 64'h5000000004000000 : _GEN_41; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_43 = 9'h2b == index ? 64'h300000000f15365 : _GEN_42; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_44 = 9'h2c == index ? 64'h1b00000017000000 : _GEN_43; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_45 = 9'h2d == index ? 64'h726777686e65706f : _GEN_44; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_46 = 9'h2e == index ? 64'h366176632c70756f : _GEN_45; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_47 = 9'h2f == index ? 64'h766373697200 : _GEN_46; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_48 = 9'h30 == index ? 64'h400000003000000 : _GEN_47; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_49 = 9'h31 == index ? 64'h4000000060000000 : _GEN_48; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_50 = 9'h32 == index ? 64'h400000003000000 : _GEN_49; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_51 = 9'h33 == index ? 64'h4000000073000000 : _GEN_50; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_52 = 9'h34 == index ? 64'h400000003000000 : _GEN_51; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_53 = 9'h35 == index ? 64'h40000080000000 : _GEN_52; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_54 = 9'h36 == index ? 64'h400000003000000 : _GEN_53; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_55 = 9'h37 == index ? 64'h10000008d000000 : _GEN_54; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_56 = 9'h38 == index ? 64'h400000003000000 : _GEN_55; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_57 = 9'h39 == index ? 64'h2000000098000000 : _GEN_56; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_58 = 9'h3a == index ? 64'h400000003000000 : _GEN_57; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_59 = 9'h3b == index ? 64'h757063a3000000 : _GEN_58; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_60 = 9'h3c == index ? 64'h400000003000000 : _GEN_59; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_61 = 9'h3d == index ? 64'haf000000 : _GEN_60; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_62 = 9'h3e == index ? 64'h400000003000000 : _GEN_61; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_63 = 9'h3f == index ? 64'h40000000ce000000 : _GEN_62; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_64 = 9'h40 == index ? 64'h400000003000000 : _GEN_63; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_65 = 9'h41 == index ? 64'h40000000e1000000 : _GEN_64; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_66 = 9'h42 == index ? 64'h400000003000000 : _GEN_65; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_67 = 9'h43 == index ? 64'h400000ee000000 : _GEN_66; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_68 = 9'h44 == index ? 64'h400000003000000 : _GEN_67; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_69 = 9'h45 == index ? 64'h1000000fb000000 : _GEN_68; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_70 = 9'h46 == index ? 64'h400000003000000 : _GEN_69; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_71 = 9'h47 == index ? 64'h2000000006010000 : _GEN_70; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_72 = 9'h48 == index ? 64'hb00000003000000 : _GEN_71; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_73 = 9'h49 == index ? 64'h6373697211010000 : _GEN_72; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_74 = 9'h4a == index ? 64'h393376732c76 : _GEN_73; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_75 = 9'h4b == index ? 64'h400000003000000 : _GEN_74; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_76 = 9'h4c == index ? 64'h10000001a010000 : _GEN_75; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_77 = 9'h4d == index ? 64'h400000003000000 : _GEN_76; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_78 = 9'h4e == index ? 64'h2b010000 : _GEN_77; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_79 = 9'h4f == index ? 64'hb00000003000000 : _GEN_78; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_80 = 9'h50 == index ? 64'h343676722f010000 : _GEN_79; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_81 = 9'h51 == index ? 64'h636466616d69 : _GEN_80; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_82 = 9'h52 == index ? 64'h500000003000000 : _GEN_81; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_83 = 9'h53 == index ? 64'h79616b6f39010000 : _GEN_82; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_84 = 9'h54 == index ? 64'h300000000000000 : _GEN_83; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_85 = 9'h55 == index ? 64'h3d00000004000000 : _GEN_84; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_86 = 9'h56 == index ? 64'h300000040420f00 : _GEN_85; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_87 = 9'h57 == index ? 64'h4001000000000000 : _GEN_86; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_88 = 9'h58 == index ? 64'h65746e6901000000 : _GEN_87; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_89 = 9'h59 == index ? 64'h6f632d7470757272 : _GEN_88; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_90 = 9'h5a == index ? 64'h72656c6c6f72746e : _GEN_89; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_91 = 9'h5b == index ? 64'h300000000000000 : _GEN_90; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_92 = 9'h5c == index ? 64'h4a01000004000000 : _GEN_91; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_93 = 9'h5d == index ? 64'h300000001000000 : _GEN_92; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_94 = 9'h5e == index ? 64'h1b0000000f000000 : _GEN_93; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_95 = 9'h5f == index ? 64'h70632c7663736972 : _GEN_94; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_96 = 9'h60 == index ? 64'h63746e692d75 : _GEN_95; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_97 = 9'h61 == index ? 64'h3000000 : _GEN_96; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_98 = 9'h62 == index ? 64'h30000005b010000 : _GEN_97; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_99 = 9'h63 == index ? 64'h7001000004000000 : _GEN_98; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_100 = 9'h64 == index ? 64'h200000002000000 : _GEN_99; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_101 = 9'h65 == index ? 64'h200000002000000 : _GEN_100; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_102 = 9'h66 == index ? 64'h6f6d656d01000000 : _GEN_101; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_103 = 9'h67 == index ? 64'h3030303038407972 : _GEN_102; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_104 = 9'h68 == index ? 64'h300000000303030 : _GEN_103; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_105 = 9'h69 == index ? 64'ha300000007000000 : _GEN_104; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_106 = 9'h6a == index ? 64'h79726f6d656d : _GEN_105; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_107 = 9'h6b == index ? 64'h800000003000000 : _GEN_106; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_108 = 9'h6c == index ? 64'h802b010000 : _GEN_107; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_109 = 9'h6d == index ? 64'h300000000000080 : _GEN_108; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_110 = 9'h6e == index ? 64'h7001000004000000 : _GEN_109; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_111 = 9'h6f == index ? 64'h200000001000000 : _GEN_110; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_112 = 9'h70 == index ? 64'h636f7301000000 : _GEN_111; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_113 = 9'h71 == index ? 64'h400000003000000 : _GEN_112; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_114 = 9'h72 == index ? 64'h100000000000000 : _GEN_113; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_115 = 9'h73 == index ? 64'h400000003000000 : _GEN_114; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_116 = 9'h74 == index ? 64'h10000000f000000 : _GEN_115; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_117 = 9'h75 == index ? 64'h1c00000003000000 : _GEN_116; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_118 = 9'h76 == index ? 64'h2c766a7a1b000000 : _GEN_117; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_119 = 9'h77 == index ? 64'h7069687372617473 : _GEN_118; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_120 = 9'h78 == index ? 64'h6d697300636f732d : _GEN_119; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_121 = 9'h79 == index ? 64'h7375622d656c70 : _GEN_120; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_122 = 9'h7a == index ? 64'h3000000 : _GEN_121; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_123 = 9'h7b == index ? 64'h100000078010000 : _GEN_122; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_124 = 9'h7c == index ? 64'h303240746e696c63 : _GEN_123; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_125 = 9'h7d == index ? 64'h3030303030 : _GEN_124; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_126 = 9'h7e == index ? 64'hd00000003000000 : _GEN_125; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_127 = 9'h7f == index ? 64'h637369721b000000 : _GEN_126; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_128 = 9'h80 == index ? 64'h30746e696c632c76 : _GEN_127; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_129 = 9'h81 == index ? 64'h300000000000000 : _GEN_128; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_130 = 9'h82 == index ? 64'h7f01000010000000 : _GEN_129; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_131 = 9'h83 == index ? 64'h300000002000000 : _GEN_130; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_132 = 9'h84 == index ? 64'h700000002000000 : _GEN_131; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_133 = 9'h85 == index ? 64'h800000003000000 : _GEN_132; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_134 = 9'h86 == index ? 64'h22b010000 : _GEN_133; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_135 = 9'h87 == index ? 64'h300000000000100 : _GEN_134; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_136 = 9'h88 == index ? 64'h9301000008000000 : _GEN_135; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_137 = 9'h89 == index ? 64'h6c6f72746e6f63 : _GEN_136; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_138 = 9'h8a == index ? 64'h100000002000000 : _GEN_137; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_139 = 9'h8b == index ? 64'h65642d726f727265 : _GEN_138; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_140 = 9'h8c == index ? 64'h3030334065636976 : _GEN_139; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_141 = 9'h8d == index ? 64'h300000000000030 : _GEN_140; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_142 = 9'h8e == index ? 64'h1b0000000e000000 : _GEN_141; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_143 = 9'h8f == index ? 64'h652c657669666973 : _GEN_142; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_144 = 9'h90 == index ? 64'h30726f7272 : _GEN_143; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_145 = 9'h91 == index ? 64'h800000003000000 : _GEN_144; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_146 = 9'h92 == index ? 64'h3000002b010000 : _GEN_145; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_147 = 9'h93 == index ? 64'h200000000100000 : _GEN_146; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_148 = 9'h94 == index ? 64'h65746e6901000000 : _GEN_147; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_149 = 9'h95 == index ? 64'h6f632d7470757272 : _GEN_148; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_150 = 9'h96 == index ? 64'h72656c6c6f72746e : _GEN_149; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_151 = 9'h97 == index ? 64'h3030303030306340 : _GEN_150; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_152 = 9'h98 == index ? 64'h300000000000000 : _GEN_151; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_153 = 9'h99 == index ? 64'h4a01000004000000 : _GEN_152; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_154 = 9'h9a == index ? 64'h300000001000000 : _GEN_153; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_155 = 9'h9b == index ? 64'h1b0000000c000000 : _GEN_154; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_156 = 9'h9c == index ? 64'h6c702c7663736972 : _GEN_155; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_157 = 9'h9d == index ? 64'h300000000306369 : _GEN_156; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_158 = 9'h9e == index ? 64'h5b01000000000000 : _GEN_157; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_159 = 9'h9f == index ? 64'h1000000003000000 : _GEN_158; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_160 = 9'ha0 == index ? 64'h20000007f010000 : _GEN_159; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_161 = 9'ha1 == index ? 64'h20000000b000000 : _GEN_160; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_162 = 9'ha2 == index ? 64'h300000009000000 : _GEN_161; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_163 = 9'ha3 == index ? 64'h2b01000008000000 : _GEN_162; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_164 = 9'ha4 == index ? 64'h40000000c : _GEN_163; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_165 = 9'ha5 == index ? 64'h800000003000000 : _GEN_164; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_166 = 9'ha6 == index ? 64'h746e6f6393010000 : _GEN_165; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_167 = 9'ha7 == index ? 64'h3000000006c6f72 : _GEN_166; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_168 = 9'ha8 == index ? 64'h9d01000004000000 : _GEN_167; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_169 = 9'ha9 == index ? 64'h300000001000000 : _GEN_168; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_170 = 9'haa == index ? 64'hb001000004000000 : _GEN_169; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_171 = 9'hab == index ? 64'h300000001000000 : _GEN_170; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_172 = 9'hac == index ? 64'h7001000004000000 : _GEN_171; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_173 = 9'had == index ? 64'h200000004000000 : _GEN_172; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_174 = 9'hae == index ? 64'h6967616d01000000 : _GEN_173; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_175 = 9'haf == index ? 64'h300000000304063 : _GEN_174; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_176 = 9'hb0 == index ? 64'h1b00000018000000 : _GEN_175; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_177 = 9'hb1 == index ? 64'h726174732c766a7a : _GEN_176; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_178 = 9'hb2 == index ? 64'h7a75662c70696873 : _GEN_177; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_179 = 9'hb3 == index ? 64'h636967616d2d7a : _GEN_178; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_180 = 9'hb4 == index ? 64'h800000003000000 : _GEN_179; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_181 = 9'hb5 == index ? 64'h2b010000 : _GEN_180; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_182 = 9'hb6 == index ? 64'h300000000100000 : _GEN_181; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_183 = 9'hb7 == index ? 64'h9301000008000000 : _GEN_182; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_184 = 9'hb8 == index ? 64'h6c6f72746e6f63 : _GEN_183; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_185 = 9'hb9 == index ? 64'h100000002000000 : _GEN_184; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_186 = 9'hba == index ? 64'h30303031406d6f72 : _GEN_185; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_187 = 9'hbb == index ? 64'h300000000000030 : _GEN_186; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_188 = 9'hbc == index ? 64'h1b0000000c000000 : _GEN_187; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_189 = 9'hbd == index ? 64'h722c657669666973 : _GEN_188; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_190 = 9'hbe == index ? 64'h300000000306d6f : _GEN_189; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_191 = 9'hbf == index ? 64'h2b01000008000000 : _GEN_190; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_192 = 9'hc0 == index ? 64'h10000000100 : _GEN_191; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_193 = 9'hc1 == index ? 64'h400000003000000 : _GEN_192; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_194 = 9'hc2 == index ? 64'h6d656d93010000 : _GEN_193; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_195 = 9'hc3 == index ? 64'h100000002000000 : _GEN_194; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_196 = 9'hc4 == index ? 64'h30303032406d6f72 : _GEN_195; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_197 = 9'hc5 == index ? 64'h300000000000030 : _GEN_196; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_198 = 9'hc6 == index ? 64'h1b00000010000000 : _GEN_197; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_199 = 9'hc7 == index ? 64'h6d2c657669666973 : _GEN_198; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_200 = 9'hc8 == index ? 64'h306d6f726b7361 : _GEN_199; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_201 = 9'hc9 == index ? 64'h800000003000000 : _GEN_200; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_202 = 9'hca == index ? 64'h2002b010000 : _GEN_201; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_203 = 9'hcb == index ? 64'h300000000200000 : _GEN_202; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_204 = 9'hcc == index ? 64'h9301000004000000 : _GEN_203; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_205 = 9'hcd == index ? 64'h2000000006d656d : _GEN_204; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_206 = 9'hce == index ? 64'h6972657301000000 : _GEN_205; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_207 = 9'hcf == index ? 64'h3030303436406c61 : _GEN_206; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_208 = 9'hd0 == index ? 64'h300000000303030 : _GEN_207; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_209 = 9'hd1 == index ? 64'hbb01000004000000 : _GEN_208; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_210 = 9'hd2 == index ? 64'h300000003000000 : _GEN_209; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_211 = 9'hd3 == index ? 64'h1b0000000d000000 : _GEN_210; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_212 = 9'hd4 == index ? 64'h752c657669666973 : _GEN_211; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_213 = 9'hd5 == index ? 64'h30747261 : _GEN_212; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_214 = 9'hd6 == index ? 64'h400000003000000 : _GEN_213; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_215 = 9'hd7 == index ? 64'h4000000c2010000 : _GEN_214; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_216 = 9'hd8 == index ? 64'h400000003000000 : _GEN_215; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_217 = 9'hd9 == index ? 64'h1000000d3010000 : _GEN_216; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_218 = 9'hda == index ? 64'h800000003000000 : _GEN_217; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_219 = 9'hdb == index ? 64'h642b010000 : _GEN_218; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_220 = 9'hdc == index ? 64'h300000000100000 : _GEN_219; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_221 = 9'hdd == index ? 64'h9301000008000000 : _GEN_220; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_222 = 9'hde == index ? 64'h6c6f72746e6f63 : _GEN_221; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_223 = 9'hdf == index ? 64'h100000002000000 : _GEN_222; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_224 = 9'he0 == index ? 64'h6574737973627573 : _GEN_223; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_225 = 9'he1 == index ? 64'h635f737562705f6d : _GEN_224; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_226 = 9'he2 == index ? 64'h6b636f6c : _GEN_225; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_227 = 9'he3 == index ? 64'h400000003000000 : _GEN_226; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_228 = 9'he4 == index ? 64'hde010000 : _GEN_227; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_229 = 9'he5 == index ? 64'h400000003000000 : _GEN_228; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_230 = 9'he6 == index ? 64'he1f50550000000 : _GEN_229; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_231 = 9'he7 == index ? 64'h1500000003000000 : _GEN_230; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_232 = 9'he8 == index ? 64'h73627573eb010000 : _GEN_231; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_233 = 9'he9 == index ? 64'h62705f6d65747379 : _GEN_232; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_234 = 9'hea == index ? 64'h6b636f6c635f7375 : _GEN_233; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_235 = 9'heb == index ? 64'h300000000000000 : _GEN_234; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_236 = 9'hec == index ? 64'h1b0000000c000000 : _GEN_235; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_237 = 9'hed == index ? 64'h6c632d6465786966 : _GEN_236; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_238 = 9'hee == index ? 64'h3000000006b636f : _GEN_237; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_239 = 9'hef == index ? 64'h7001000004000000 : _GEN_238; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_240 = 9'hf0 == index ? 64'h200000003000000 : _GEN_239; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_241 = 9'hf1 == index ? 64'h200000002000000 : _GEN_240; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_242 = 9'hf2 == index ? 64'h6464612309000000 : _GEN_241; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_243 = 9'hf3 == index ? 64'h6c65632d73736572 : _GEN_242; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_244 = 9'hf4 == index ? 64'h657a69732300736c : _GEN_243; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_245 = 9'hf5 == index ? 64'h6300736c6c65632d : _GEN_244; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_246 = 9'hf6 == index ? 64'h6c62697461706d6f : _GEN_245; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_247 = 9'hf7 == index ? 64'h6c65646f6d0065 : _GEN_246; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_248 = 9'hf8 == index ? 64'h306c6169726573 : _GEN_247; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_249 = 9'hf9 == index ? 64'h73677261746f6f62 : _GEN_248; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_250 = 9'hfa == index ? 64'h736162656d697400 : _GEN_249; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_251 = 9'hfb == index ? 64'h6575716572662d65 : _GEN_250; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_252 = 9'hfc == index ? 64'h636f6c630079636e : _GEN_251; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_253 = 9'hfd == index ? 64'h6575716572662d6b : _GEN_252; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_254 = 9'hfe == index ? 64'h61632d640079636e : _GEN_253; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_255 = 9'hff == index ? 64'h636f6c622d656863 : _GEN_254; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_256 = 9'h100 == index ? 64'h6400657a69732d6b : _GEN_255; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_257 = 9'h101 == index ? 64'h732d65686361632d : _GEN_256; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_258 = 9'h102 == index ? 64'h61632d6400737465 : _GEN_257; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_259 = 9'h103 == index ? 64'h657a69732d656863 : _GEN_258; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_260 = 9'h104 == index ? 64'h732d626c742d6400 : _GEN_259; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_261 = 9'h105 == index ? 64'h6c742d6400737465 : _GEN_260; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_262 = 9'h106 == index ? 64'h6400657a69732d62 : _GEN_261; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_263 = 9'h107 == index ? 64'h79745f6563697665 : _GEN_262; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_264 = 9'h108 == index ? 64'h7764726168006570 : _GEN_263; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_265 = 9'h109 == index ? 64'h636578652d657261 : _GEN_264; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_266 = 9'h10a == index ? 64'h6f706b616572622d : _GEN_265; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_267 = 9'h10b == index ? 64'h6e756f632d746e69 : _GEN_266; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_268 = 9'h10c == index ? 64'h686361632d690074 : _GEN_267; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_269 = 9'h10d == index ? 64'h2d6b636f6c622d65 : _GEN_268; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_270 = 9'h10e == index ? 64'h632d6900657a6973 : _GEN_269; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_271 = 9'h10f == index ? 64'h7465732d65686361 : _GEN_270; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_272 = 9'h110 == index ? 64'h686361632d690073 : _GEN_271; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_273 = 9'h111 == index ? 64'h6900657a69732d65 : _GEN_272; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_274 = 9'h112 == index ? 64'h7465732d626c742d : _GEN_273; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_275 = 9'h113 == index ? 64'h2d626c742d690073 : _GEN_274; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_276 = 9'h114 == index ? 64'h756d6d00657a6973 : _GEN_275; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_277 = 9'h115 == index ? 64'h656e00657079742d : _GEN_276; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_278 = 9'h116 == index ? 64'h6c6576656c2d7478 : _GEN_277; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_279 = 9'h117 == index ? 64'h720065686361632d : _GEN_278; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_280 = 9'h118 == index ? 64'h7663736972006765 : _GEN_279; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_281 = 9'h119 == index ? 64'h617473006173692c : _GEN_280; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_282 = 9'h11a == index ? 64'h2d626c7400737574 : _GEN_281; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_283 = 9'h11b == index ? 64'h69230074696c7073 : _GEN_282; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_284 = 9'h11c == index ? 64'h747075727265746e : _GEN_283; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_285 = 9'h11d == index ? 64'h6900736c6c65632d : _GEN_284; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_286 = 9'h11e == index ? 64'h747075727265746e : _GEN_285; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_287 = 9'h11f == index ? 64'h6c6f72746e6f632d : _GEN_286; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_288 = 9'h120 == index ? 64'h6e6168700072656c : _GEN_287; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_289 = 9'h121 == index ? 64'h676e617200656c64 : _GEN_288; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_290 = 9'h122 == index ? 64'h7265746e69007365 : _GEN_289; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_291 = 9'h123 == index ? 64'h78652d7374707572 : _GEN_290; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_292 = 9'h124 == index ? 64'h72006465646e6574 : _GEN_291; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_293 = 9'h125 == index ? 64'h73656d616e2d6765 : _GEN_292; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_294 = 9'h126 == index ? 64'h6d2c766373697200 : _GEN_293; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_295 = 9'h127 == index ? 64'h726f6972702d7861 : _GEN_294; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_296 = 9'h128 == index ? 64'h6373697200797469 : _GEN_295; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_297 = 9'h129 == index ? 64'h63007665646e2c76 : _GEN_296; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_298 = 9'h12a == index ? 64'h6e6900736b636f6c : _GEN_297; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_299 = 9'h12b == index ? 64'h2d74707572726574 : _GEN_298; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_300 = 9'h12c == index ? 64'h6900746e65726170 : _GEN_299; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_301 = 9'h12d == index ? 64'h747075727265746e : _GEN_300; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_302 = 9'h12e == index ? 64'h6b636f6c63230073 : _GEN_301; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_303 = 9'h12f == index ? 64'h6300736c6c65632d : _GEN_302; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_304 = 9'h130 == index ? 64'h74756f2d6b636f6c : _GEN_303; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_305 = 9'h131 == index ? 64'h656d616e2d747570 : _GEN_304; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_306 = 9'h132 == index ? 64'h73 : _GEN_305; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_307 = 9'h133 == index ? 64'h0 : _GEN_306; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_308 = 9'h134 == index ? 64'h0 : _GEN_307; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_309 = 9'h135 == index ? 64'h0 : _GEN_308; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_310 = 9'h136 == index ? 64'h0 : _GEN_309; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_311 = 9'h137 == index ? 64'h0 : _GEN_310; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_312 = 9'h138 == index ? 64'h0 : _GEN_311; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_313 = 9'h139 == index ? 64'h0 : _GEN_312; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_314 = 9'h13a == index ? 64'h0 : _GEN_313; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_315 = 9'h13b == index ? 64'h0 : _GEN_314; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_316 = 9'h13c == index ? 64'h0 : _GEN_315; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_317 = 9'h13d == index ? 64'h0 : _GEN_316; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_318 = 9'h13e == index ? 64'h0 : _GEN_317; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_319 = 9'h13f == index ? 64'h0 : _GEN_318; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_320 = 9'h140 == index ? 64'h0 : _GEN_319; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_321 = 9'h141 == index ? 64'h0 : _GEN_320; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_322 = 9'h142 == index ? 64'h0 : _GEN_321; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_323 = 9'h143 == index ? 64'h0 : _GEN_322; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_324 = 9'h144 == index ? 64'h0 : _GEN_323; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_325 = 9'h145 == index ? 64'h0 : _GEN_324; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_326 = 9'h146 == index ? 64'h0 : _GEN_325; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_327 = 9'h147 == index ? 64'h0 : _GEN_326; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_328 = 9'h148 == index ? 64'h0 : _GEN_327; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_329 = 9'h149 == index ? 64'h0 : _GEN_328; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_330 = 9'h14a == index ? 64'h0 : _GEN_329; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_331 = 9'h14b == index ? 64'h0 : _GEN_330; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_332 = 9'h14c == index ? 64'h0 : _GEN_331; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_333 = 9'h14d == index ? 64'h0 : _GEN_332; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_334 = 9'h14e == index ? 64'h0 : _GEN_333; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_335 = 9'h14f == index ? 64'h0 : _GEN_334; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_336 = 9'h150 == index ? 64'h0 : _GEN_335; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_337 = 9'h151 == index ? 64'h0 : _GEN_336; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_338 = 9'h152 == index ? 64'h0 : _GEN_337; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_339 = 9'h153 == index ? 64'h0 : _GEN_338; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_340 = 9'h154 == index ? 64'h0 : _GEN_339; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_341 = 9'h155 == index ? 64'h0 : _GEN_340; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_342 = 9'h156 == index ? 64'h0 : _GEN_341; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_343 = 9'h157 == index ? 64'h0 : _GEN_342; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_344 = 9'h158 == index ? 64'h0 : _GEN_343; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_345 = 9'h159 == index ? 64'h0 : _GEN_344; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_346 = 9'h15a == index ? 64'h0 : _GEN_345; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_347 = 9'h15b == index ? 64'h0 : _GEN_346; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_348 = 9'h15c == index ? 64'h0 : _GEN_347; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_349 = 9'h15d == index ? 64'h0 : _GEN_348; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_350 = 9'h15e == index ? 64'h0 : _GEN_349; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_351 = 9'h15f == index ? 64'h0 : _GEN_350; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_352 = 9'h160 == index ? 64'h0 : _GEN_351; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_353 = 9'h161 == index ? 64'h0 : _GEN_352; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_354 = 9'h162 == index ? 64'h0 : _GEN_353; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_355 = 9'h163 == index ? 64'h0 : _GEN_354; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_356 = 9'h164 == index ? 64'h0 : _GEN_355; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_357 = 9'h165 == index ? 64'h0 : _GEN_356; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_358 = 9'h166 == index ? 64'h0 : _GEN_357; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_359 = 9'h167 == index ? 64'h0 : _GEN_358; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_360 = 9'h168 == index ? 64'h0 : _GEN_359; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_361 = 9'h169 == index ? 64'h0 : _GEN_360; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_362 = 9'h16a == index ? 64'h0 : _GEN_361; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_363 = 9'h16b == index ? 64'h0 : _GEN_362; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_364 = 9'h16c == index ? 64'h0 : _GEN_363; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_365 = 9'h16d == index ? 64'h0 : _GEN_364; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_366 = 9'h16e == index ? 64'h0 : _GEN_365; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_367 = 9'h16f == index ? 64'h0 : _GEN_366; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_368 = 9'h170 == index ? 64'h0 : _GEN_367; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_369 = 9'h171 == index ? 64'h0 : _GEN_368; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_370 = 9'h172 == index ? 64'h0 : _GEN_369; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_371 = 9'h173 == index ? 64'h0 : _GEN_370; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_372 = 9'h174 == index ? 64'h0 : _GEN_371; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_373 = 9'h175 == index ? 64'h0 : _GEN_372; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_374 = 9'h176 == index ? 64'h0 : _GEN_373; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_375 = 9'h177 == index ? 64'h0 : _GEN_374; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_376 = 9'h178 == index ? 64'h0 : _GEN_375; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_377 = 9'h179 == index ? 64'h0 : _GEN_376; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_378 = 9'h17a == index ? 64'h0 : _GEN_377; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_379 = 9'h17b == index ? 64'h0 : _GEN_378; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_380 = 9'h17c == index ? 64'h0 : _GEN_379; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_381 = 9'h17d == index ? 64'h0 : _GEN_380; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_382 = 9'h17e == index ? 64'h0 : _GEN_381; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_383 = 9'h17f == index ? 64'h0 : _GEN_382; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_384 = 9'h180 == index ? 64'h0 : _GEN_383; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_385 = 9'h181 == index ? 64'h0 : _GEN_384; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_386 = 9'h182 == index ? 64'h0 : _GEN_385; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_387 = 9'h183 == index ? 64'h0 : _GEN_386; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_388 = 9'h184 == index ? 64'h0 : _GEN_387; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_389 = 9'h185 == index ? 64'h0 : _GEN_388; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_390 = 9'h186 == index ? 64'h0 : _GEN_389; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_391 = 9'h187 == index ? 64'h0 : _GEN_390; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_392 = 9'h188 == index ? 64'h0 : _GEN_391; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_393 = 9'h189 == index ? 64'h0 : _GEN_392; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_394 = 9'h18a == index ? 64'h0 : _GEN_393; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_395 = 9'h18b == index ? 64'h0 : _GEN_394; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_396 = 9'h18c == index ? 64'h0 : _GEN_395; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_397 = 9'h18d == index ? 64'h0 : _GEN_396; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_398 = 9'h18e == index ? 64'h0 : _GEN_397; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_399 = 9'h18f == index ? 64'h0 : _GEN_398; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_400 = 9'h190 == index ? 64'h0 : _GEN_399; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_401 = 9'h191 == index ? 64'h0 : _GEN_400; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_402 = 9'h192 == index ? 64'h0 : _GEN_401; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_403 = 9'h193 == index ? 64'h0 : _GEN_402; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_404 = 9'h194 == index ? 64'h0 : _GEN_403; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_405 = 9'h195 == index ? 64'h0 : _GEN_404; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_406 = 9'h196 == index ? 64'h0 : _GEN_405; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_407 = 9'h197 == index ? 64'h0 : _GEN_406; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_408 = 9'h198 == index ? 64'h0 : _GEN_407; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_409 = 9'h199 == index ? 64'h0 : _GEN_408; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_410 = 9'h19a == index ? 64'h0 : _GEN_409; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_411 = 9'h19b == index ? 64'h0 : _GEN_410; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_412 = 9'h19c == index ? 64'h0 : _GEN_411; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_413 = 9'h19d == index ? 64'h0 : _GEN_412; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_414 = 9'h19e == index ? 64'h0 : _GEN_413; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_415 = 9'h19f == index ? 64'h0 : _GEN_414; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_416 = 9'h1a0 == index ? 64'h0 : _GEN_415; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_417 = 9'h1a1 == index ? 64'h0 : _GEN_416; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_418 = 9'h1a2 == index ? 64'h0 : _GEN_417; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_419 = 9'h1a3 == index ? 64'h0 : _GEN_418; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_420 = 9'h1a4 == index ? 64'h0 : _GEN_419; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_421 = 9'h1a5 == index ? 64'h0 : _GEN_420; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_422 = 9'h1a6 == index ? 64'h0 : _GEN_421; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_423 = 9'h1a7 == index ? 64'h0 : _GEN_422; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_424 = 9'h1a8 == index ? 64'h0 : _GEN_423; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_425 = 9'h1a9 == index ? 64'h0 : _GEN_424; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_426 = 9'h1aa == index ? 64'h0 : _GEN_425; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_427 = 9'h1ab == index ? 64'h0 : _GEN_426; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_428 = 9'h1ac == index ? 64'h0 : _GEN_427; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_429 = 9'h1ad == index ? 64'h0 : _GEN_428; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_430 = 9'h1ae == index ? 64'h0 : _GEN_429; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_431 = 9'h1af == index ? 64'h0 : _GEN_430; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_432 = 9'h1b0 == index ? 64'h0 : _GEN_431; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_433 = 9'h1b1 == index ? 64'h0 : _GEN_432; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_434 = 9'h1b2 == index ? 64'h0 : _GEN_433; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_435 = 9'h1b3 == index ? 64'h0 : _GEN_434; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_436 = 9'h1b4 == index ? 64'h0 : _GEN_435; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_437 = 9'h1b5 == index ? 64'h0 : _GEN_436; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_438 = 9'h1b6 == index ? 64'h0 : _GEN_437; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_439 = 9'h1b7 == index ? 64'h0 : _GEN_438; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_440 = 9'h1b8 == index ? 64'h0 : _GEN_439; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_441 = 9'h1b9 == index ? 64'h0 : _GEN_440; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_442 = 9'h1ba == index ? 64'h0 : _GEN_441; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_443 = 9'h1bb == index ? 64'h0 : _GEN_442; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_444 = 9'h1bc == index ? 64'h0 : _GEN_443; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_445 = 9'h1bd == index ? 64'h0 : _GEN_444; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_446 = 9'h1be == index ? 64'h0 : _GEN_445; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_447 = 9'h1bf == index ? 64'h0 : _GEN_446; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_448 = 9'h1c0 == index ? 64'h0 : _GEN_447; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_449 = 9'h1c1 == index ? 64'h0 : _GEN_448; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_450 = 9'h1c2 == index ? 64'h0 : _GEN_449; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_451 = 9'h1c3 == index ? 64'h0 : _GEN_450; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_452 = 9'h1c4 == index ? 64'h0 : _GEN_451; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_453 = 9'h1c5 == index ? 64'h0 : _GEN_452; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_454 = 9'h1c6 == index ? 64'h0 : _GEN_453; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_455 = 9'h1c7 == index ? 64'h0 : _GEN_454; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_456 = 9'h1c8 == index ? 64'h0 : _GEN_455; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_457 = 9'h1c9 == index ? 64'h0 : _GEN_456; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_458 = 9'h1ca == index ? 64'h0 : _GEN_457; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_459 = 9'h1cb == index ? 64'h0 : _GEN_458; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_460 = 9'h1cc == index ? 64'h0 : _GEN_459; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_461 = 9'h1cd == index ? 64'h0 : _GEN_460; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_462 = 9'h1ce == index ? 64'h0 : _GEN_461; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_463 = 9'h1cf == index ? 64'h0 : _GEN_462; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_464 = 9'h1d0 == index ? 64'h0 : _GEN_463; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_465 = 9'h1d1 == index ? 64'h0 : _GEN_464; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_466 = 9'h1d2 == index ? 64'h0 : _GEN_465; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_467 = 9'h1d3 == index ? 64'h0 : _GEN_466; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_468 = 9'h1d4 == index ? 64'h0 : _GEN_467; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_469 = 9'h1d5 == index ? 64'h0 : _GEN_468; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_470 = 9'h1d6 == index ? 64'h0 : _GEN_469; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_471 = 9'h1d7 == index ? 64'h0 : _GEN_470; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_472 = 9'h1d8 == index ? 64'h0 : _GEN_471; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_473 = 9'h1d9 == index ? 64'h0 : _GEN_472; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_474 = 9'h1da == index ? 64'h0 : _GEN_473; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_475 = 9'h1db == index ? 64'h0 : _GEN_474; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_476 = 9'h1dc == index ? 64'h0 : _GEN_475; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_477 = 9'h1dd == index ? 64'h0 : _GEN_476; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_478 = 9'h1de == index ? 64'h0 : _GEN_477; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_479 = 9'h1df == index ? 64'h0 : _GEN_478; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_480 = 9'h1e0 == index ? 64'h0 : _GEN_479; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_481 = 9'h1e1 == index ? 64'h0 : _GEN_480; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_482 = 9'h1e2 == index ? 64'h0 : _GEN_481; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_483 = 9'h1e3 == index ? 64'h0 : _GEN_482; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_484 = 9'h1e4 == index ? 64'h0 : _GEN_483; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_485 = 9'h1e5 == index ? 64'h0 : _GEN_484; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_486 = 9'h1e6 == index ? 64'h0 : _GEN_485; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_487 = 9'h1e7 == index ? 64'h0 : _GEN_486; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_488 = 9'h1e8 == index ? 64'h0 : _GEN_487; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_489 = 9'h1e9 == index ? 64'h0 : _GEN_488; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_490 = 9'h1ea == index ? 64'h0 : _GEN_489; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_491 = 9'h1eb == index ? 64'h0 : _GEN_490; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_492 = 9'h1ec == index ? 64'h0 : _GEN_491; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_493 = 9'h1ed == index ? 64'h0 : _GEN_492; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_494 = 9'h1ee == index ? 64'h0 : _GEN_493; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_495 = 9'h1ef == index ? 64'h0 : _GEN_494; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_496 = 9'h1f0 == index ? 64'h0 : _GEN_495; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_497 = 9'h1f1 == index ? 64'h0 : _GEN_496; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_498 = 9'h1f2 == index ? 64'h0 : _GEN_497; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_499 = 9'h1f3 == index ? 64'h0 : _GEN_498; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_500 = 9'h1f4 == index ? 64'h0 : _GEN_499; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_501 = 9'h1f5 == index ? 64'h0 : _GEN_500; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_502 = 9'h1f6 == index ? 64'h0 : _GEN_501; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_503 = 9'h1f7 == index ? 64'h0 : _GEN_502; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_504 = 9'h1f8 == index ? 64'h0 : _GEN_503; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_505 = 9'h1f9 == index ? 64'h0 : _GEN_504; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_506 = 9'h1fa == index ? 64'h0 : _GEN_505; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_507 = 9'h1fb == index ? 64'h0 : _GEN_506; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_508 = 9'h1fc == index ? 64'h0 : _GEN_507; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_509 = 9'h1fd == index ? 64'h0 : _GEN_508; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_510 = 9'h1fe == index ? 64'h0 : _GEN_509; // @[BootROM.scala 51:{47,47}]
  wire [63:0] _GEN_511 = 9'h1ff == index ? 64'h0 : _GEN_510; // @[BootROM.scala 51:{47,47}]
  wire [29:0] TLROM_covSum;
  assign auto_in_a_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_in_d_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_in_d_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_in_d_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_in_d_bits_data = |high ? 64'h0 : _GEN_511; // @[BootROM.scala 51:47]
  assign TLROM_covSum = 30'h0;
  assign io_covSum = TLROM_covSum;
endmodule
module ClockSinkDomain_1(
  output        auto_bootrom_in_a_ready,
  input         auto_bootrom_in_a_valid,
  input  [1:0]  auto_bootrom_in_a_bits_size,
  input  [10:0] auto_bootrom_in_a_bits_source,
  input  [16:0] auto_bootrom_in_a_bits_address,
  input         auto_bootrom_in_d_ready,
  output        auto_bootrom_in_d_valid,
  output [1:0]  auto_bootrom_in_d_bits_size,
  output [10:0] auto_bootrom_in_d_bits_source,
  output [63:0] auto_bootrom_in_d_bits_data,
  output [29:0] io_covSum
);
  wire  bootrom_auto_in_a_ready; // @[BootROM.scala 81:17]
  wire  bootrom_auto_in_a_valid; // @[BootROM.scala 81:17]
  wire [1:0] bootrom_auto_in_a_bits_size; // @[BootROM.scala 81:17]
  wire [10:0] bootrom_auto_in_a_bits_source; // @[BootROM.scala 81:17]
  wire [16:0] bootrom_auto_in_a_bits_address; // @[BootROM.scala 81:17]
  wire  bootrom_auto_in_d_ready; // @[BootROM.scala 81:17]
  wire  bootrom_auto_in_d_valid; // @[BootROM.scala 81:17]
  wire [1:0] bootrom_auto_in_d_bits_size; // @[BootROM.scala 81:17]
  wire [10:0] bootrom_auto_in_d_bits_source; // @[BootROM.scala 81:17]
  wire [63:0] bootrom_auto_in_d_bits_data; // @[BootROM.scala 81:17]
  wire [29:0] bootrom_io_covSum; // @[BootROM.scala 81:17]
  wire [29:0] ClockSinkDomain_1_covSum;
  wire [29:0] bootrom_sum;
  TLROM bootrom ( // @[BootROM.scala 81:17]
    .auto_in_a_ready(bootrom_auto_in_a_ready),
    .auto_in_a_valid(bootrom_auto_in_a_valid),
    .auto_in_a_bits_size(bootrom_auto_in_a_bits_size),
    .auto_in_a_bits_source(bootrom_auto_in_a_bits_source),
    .auto_in_a_bits_address(bootrom_auto_in_a_bits_address),
    .auto_in_d_ready(bootrom_auto_in_d_ready),
    .auto_in_d_valid(bootrom_auto_in_d_valid),
    .auto_in_d_bits_size(bootrom_auto_in_d_bits_size),
    .auto_in_d_bits_source(bootrom_auto_in_d_bits_source),
    .auto_in_d_bits_data(bootrom_auto_in_d_bits_data),
    .io_covSum(bootrom_io_covSum)
  );
  assign auto_bootrom_in_a_ready = bootrom_auto_in_a_ready; // @[LazyModule.scala 309:16]
  assign auto_bootrom_in_d_valid = bootrom_auto_in_d_valid; // @[LazyModule.scala 309:16]
  assign auto_bootrom_in_d_bits_size = bootrom_auto_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_bootrom_in_d_bits_source = bootrom_auto_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign auto_bootrom_in_d_bits_data = bootrom_auto_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign bootrom_auto_in_a_valid = auto_bootrom_in_a_valid; // @[LazyModule.scala 309:16]
  assign bootrom_auto_in_a_bits_size = auto_bootrom_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign bootrom_auto_in_a_bits_source = auto_bootrom_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign bootrom_auto_in_a_bits_address = auto_bootrom_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign bootrom_auto_in_d_ready = auto_bootrom_in_d_ready; // @[LazyModule.scala 309:16]
  assign ClockSinkDomain_1_covSum = 30'h0;
  assign bootrom_sum = ClockSinkDomain_1_covSum + bootrom_io_covSum;
  assign io_covSum = bootrom_sum;
endmodule
module TLMaskROM(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [1:0]  auto_in_a_bits_size,
  input  [11:0] auto_in_a_bits_source,
  input  [17:0] auto_in_a_bits_address,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [1:0]  auto_in_d_bits_size,
  output [11:0] auto_in_d_bits_source,
  output [31:0] auto_in_d_bits_data,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  rom_clock; // @[ROMGenerator.scala 27:19]
  wire [10:0] rom_address; // @[ROMGenerator.scala 27:19]
  wire  rom_oe; // @[ROMGenerator.scala 27:19]
  wire  rom_me; // @[ROMGenerator.scala 27:19]
  wire [31:0] rom_q; // @[ROMGenerator.scala 27:19]
  wire [17:0] _rom_io_address_T_1 = auto_in_a_bits_address - 18'h20000; // @[MaskROM.scala 31:54]
  reg  d_full; // @[MaskROM.scala 35:25]
  wire  in_a_ready = auto_in_d_ready | ~d_full; // @[MaskROM.scala 44:30]
  wire  _rom_io_me_T = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 50:35]
  reg [1:0] d_size; // @[MaskROM.scala 36:21]
  reg [11:0] d_source; // @[MaskROM.scala 37:23]
  reg  d_data_REG; // @[MaskROM.scala 38:45]
  reg [31:0] d_data_r; // @[Reg.scala 16:16]
  wire  _T = auto_in_d_ready & d_full; // @[Decoupled.scala 50:35]
  wire  _GEN_1 = _T ? 1'h0 : d_full; // @[MaskROM.scala 41:24 35:25 41:33]
  wire  _GEN_2 = _rom_io_me_T | _GEN_1; // @[MaskROM.scala 42:{24,33}]
  reg [1:0] TLMaskROM_covState; // @[Register tracking TLMaskROM state]
  reg  TLMaskROM_covMap [0:3]; // @[Coverage map for TLMaskROM]
  wire  TLMaskROM_covMap_read_en; // @[Coverage map for TLMaskROM]
  wire [1:0] TLMaskROM_covMap_read_addr; // @[Coverage map for TLMaskROM]
  wire  TLMaskROM_covMap_read_data; // @[Coverage map for TLMaskROM]
  wire  TLMaskROM_covMap_write_data; // @[Coverage map for TLMaskROM]
  wire [1:0] TLMaskROM_covMap_write_addr; // @[Coverage map for TLMaskROM]
  wire  TLMaskROM_covMap_write_mask; // @[Coverage map for TLMaskROM]
  wire  TLMaskROM_covMap_write_en; // @[Coverage map for TLMaskROM]
  reg [29:0] TLMaskROM_covSum; // @[Sum of coverage map]
  wire  d_data_REG_shl;
  wire [1:0] d_data_REG_pad;
  wire [1:0] d_full_shl;
  wire [1:0] d_full_pad;
  wire [1:0] TLMaskROM_xor0;
  StarshipROM rom ( // @[ROMGenerator.scala 27:19]
    .clock(rom_clock),
    .address(rom_address),
    .oe(rom_oe),
    .me(rom_me),
    .q(rom_q)
  );
  assign auto_in_a_ready = auto_in_d_ready | ~d_full; // @[MaskROM.scala 44:30]
  assign auto_in_d_valid = d_full; // @[Nodes.scala 1210:84 MaskROM.scala 43:16]
  assign auto_in_d_bits_size = d_size; // @[Edges.scala 771:17 774:15]
  assign auto_in_d_bits_source = d_source; // @[Edges.scala 771:17 775:15]
  assign auto_in_d_bits_data = d_data_REG ? rom_q : d_data_r; // @[package.scala 79:42]
  assign rom_clock = clock; // @[MaskROM.scala 30:18]
  assign rom_address = _rom_io_address_T_1[12:2]; // @[MaskROM.scala 31:72]
  assign rom_oe = 1'h1; // @[MaskROM.scala 32:15]
  assign rom_me = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 50:35]
  assign TLMaskROM_covMap_read_en = 1'h1;
  assign TLMaskROM_covMap_read_addr = TLMaskROM_covState;
  assign TLMaskROM_covMap_read_data = TLMaskROM_covMap[TLMaskROM_covMap_read_addr]; // @[Coverage map for TLMaskROM]
  assign TLMaskROM_covMap_write_data = 1'h1;
  assign TLMaskROM_covMap_write_addr = TLMaskROM_covState;
  assign TLMaskROM_covMap_write_mask = 1'h1;
  assign TLMaskROM_covMap_write_en = ~metaReset;
  assign d_data_REG_shl = d_data_REG;
  assign d_data_REG_pad = {1'h0,d_data_REG_shl};
  assign d_full_shl = {d_full, 1'h0};
  assign d_full_pad = d_full_shl;
  assign TLMaskROM_xor0 = d_data_REG_pad ^ d_full_pad;
  assign io_covSum = TLMaskROM_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[MaskROM.scala 35:25]
      d_full <= 1'h0; // @[MaskROM.scala 35:25]
    end else begin
      d_full <= _GEN_2;
    end
    if (_rom_io_me_T) begin // @[MaskROM.scala 46:24]
      d_size <= auto_in_a_bits_size; // @[MaskROM.scala 47:16]
    end
    if (_rom_io_me_T) begin // @[MaskROM.scala 46:24]
      d_source <= auto_in_a_bits_source; // @[MaskROM.scala 48:16]
    end
    d_data_REG <= in_a_ready & auto_in_a_valid; // @[Decoupled.scala 50:35]
    if (d_data_REG) begin // @[Reg.scala 17:18]
      d_data_r <= rom_q; // @[Reg.scala 17:22]
    end
    TLMaskROM_covState <= TLMaskROM_xor0;
    if (TLMaskROM_covMap_write_en & TLMaskROM_covMap_write_mask) begin
      TLMaskROM_covMap[TLMaskROM_covMap_write_addr] <= TLMaskROM_covMap_write_data; // @[Coverage map for TLMaskROM]
    end
    if (!(TLMaskROM_covMap_read_data | metaReset)) begin
      TLMaskROM_covSum <= TLMaskROM_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    TLMaskROM_covMap[initvar] = 0; //_6[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  d_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  d_size = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  d_source = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  d_data_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  d_data_r = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  TLMaskROM_covState = 0; //_5[1:0];
  _RAND_7 = {1{`RANDOM}};
  TLMaskROM_covSum = 0; //_7[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module UARTTx(
  input         clock,
  input         reset,
  input         io_en,
  output        io_in_ready,
  input         io_in_valid,
  input  [7:0]  io_in_bits,
  output        io_out,
  input  [15:0] io_div,
  input         io_nstop,
  output [29:0] io_covSum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  reg [15:0] prescaler; // @[UARTTx.scala 23:22]
  wire  pulse = prescaler == 16'h0; // @[UARTTx.scala 24:26]
  reg [3:0] counter; // @[UARTTx.scala 27:20]
  reg [8:0] shifter; // @[UARTTx.scala 28:20]
  reg  out; // @[UARTTx.scala 29:16]
  wire  plusarg_tx = |plusarg_reader_out; // @[UARTTx.scala 32:90]
  wire  busy = counter != 4'h0; // @[UARTTx.scala 34:23]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 50:35]
  wire [9:0] _shifter_T_1 = {1'h1,io_in_bits,1'h0}; // @[Cat.scala 31:58]
  wire  _counter_T = ~io_nstop; // @[UARTTx.scala 57:19]
  wire [3:0] _counter_T_2 = _counter_T ? 4'ha : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _counter_T_3 = io_nstop ? 4'hb : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _counter_T_4 = _counter_T_2 | _counter_T_3; // @[Mux.scala 27:73]
  wire [3:0] _counter_T_6 = _counter_T_4 - 4'h0; // @[UARTTx.scala 57:53]
  wire [9:0] _GEN_0 = _T & plusarg_tx ? _shifter_T_1 : {{1'd0}, shifter}; // @[UARTTx.scala 40:37 55:15 28:20]
  wire [15:0] _prescaler_T_2 = prescaler - 16'h1; // @[UARTTx.scala 61:78]
  wire [3:0] _counter_T_8 = counter - 4'h1; // @[UARTTx.scala 64:24]
  wire [8:0] _shifter_T_3 = {1'h1,shifter[8:1]}; // @[Cat.scala 31:58]
  wire [9:0] _GEN_4 = pulse & busy ? {{1'd0}, _shifter_T_3} : _GEN_0; // @[UARTTx.scala 63:24 65:13]
  wire  _GEN_5 = pulse & busy ? shifter[0] : out; // @[UARTTx.scala 29:16 63:24 66:9]
  wire [29:0] UARTTx_covSum;
  plusarg_reader #(.FORMAT("uart_tx=%d"), .DEFAULT(1), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  assign io_in_ready = io_en & ~busy; // @[UARTTx.scala 35:24]
  assign io_out = out; // @[UARTTx.scala 30:10]
  assign UARTTx_covSum = 30'h0;
  assign io_covSum = UARTTx_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[UARTTx.scala 23:22]
      prescaler <= 16'h0; // @[UARTTx.scala 23:22]
    end else if (busy) begin
      if (pulse) begin
        prescaler <= io_div;
      end else begin
        prescaler <= _prescaler_T_2;
      end
    end
    if (reset) begin // @[UARTTx.scala 27:20]
      counter <= 4'h0; // @[UARTTx.scala 27:20]
    end else if (pulse & busy) begin
      counter <= _counter_T_8;
    end else if (_T & plusarg_tx) begin
      counter <= _counter_T_6;
    end
    shifter <= _GEN_4[8:0];
    out <= reset | _GEN_5; // @[UARTTx.scala 29:{16,16}]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & ~reset) begin
          $fwrite(32'h80000002,"UART TX (%x): %c\n",io_in_bits,io_in_bits); // @[UARTTx.scala 38:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prescaler = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  shifter = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  out = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QueueCompatibility_68(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [7:0]  io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [7:0]  io_deq_bits,
  output [3:0]  io_count,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:7]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [2:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire [2:0] ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg [2:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 78:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 78:24]
  wire [2:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 312:32]
  wire [3:0] _io_count_T_1 = maybe_full & ptr_match ? 4'h8 : 4'h0; // @[Decoupled.scala 315:20]
  wire [3:0] _GEN_11 = {{1'd0}, ptr_diff}; // @[Decoupled.scala 315:62]
  reg  QueueCompatibility_68_covState; // @[Register tracking QueueCompatibility_68 state]
  reg  QueueCompatibility_68_covMap [0:1]; // @[Coverage map for QueueCompatibility_68]
  wire  QueueCompatibility_68_covMap_read_en; // @[Coverage map for QueueCompatibility_68]
  wire  QueueCompatibility_68_covMap_read_addr; // @[Coverage map for QueueCompatibility_68]
  wire  QueueCompatibility_68_covMap_read_data; // @[Coverage map for QueueCompatibility_68]
  wire  QueueCompatibility_68_covMap_write_data; // @[Coverage map for QueueCompatibility_68]
  wire  QueueCompatibility_68_covMap_write_addr; // @[Coverage map for QueueCompatibility_68]
  wire  QueueCompatibility_68_covMap_write_mask; // @[Coverage map for QueueCompatibility_68]
  wire  QueueCompatibility_68_covMap_write_en; // @[Coverage map for QueueCompatibility_68]
  reg [29:0] QueueCompatibility_68_covSum; // @[Sum of coverage map]
  wire  maybe_full_shl;
  wire  maybe_full_pad;
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_count = _io_count_T_1 | _GEN_11; // @[Decoupled.scala 315:62]
  assign QueueCompatibility_68_covMap_read_en = 1'h1;
  assign QueueCompatibility_68_covMap_read_addr = QueueCompatibility_68_covState;
  assign QueueCompatibility_68_covMap_read_data = QueueCompatibility_68_covMap[QueueCompatibility_68_covMap_read_addr]; // @[Coverage map for QueueCompatibility_68]
  assign QueueCompatibility_68_covMap_write_data = 1'h1;
  assign QueueCompatibility_68_covMap_write_addr = QueueCompatibility_68_covState;
  assign QueueCompatibility_68_covMap_write_mask = 1'h1;
  assign QueueCompatibility_68_covMap_write_en = ~metaReset;
  assign maybe_full_shl = maybe_full;
  assign maybe_full_pad = maybe_full_shl;
  assign io_covSum = QueueCompatibility_68_covSum;
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin
      enq_ptr_value <= _value_T_1;
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin
      deq_ptr_value <= _value_T_3;
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin
      maybe_full <= do_enq;
    end
    QueueCompatibility_68_covState <= maybe_full_pad;
    if (QueueCompatibility_68_covMap_write_en & QueueCompatibility_68_covMap_write_mask) begin
      QueueCompatibility_68_covMap[QueueCompatibility_68_covMap_write_addr] <= QueueCompatibility_68_covMap_write_data; // @[Coverage map for QueueCompatibility_68]
    end
    if (!(QueueCompatibility_68_covMap_read_data | metaReset)) begin
      QueueCompatibility_68_covSum <= QueueCompatibility_68_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    QueueCompatibility_68_covMap[initvar] = 0; //_5[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  QueueCompatibility_68_covState = 0; //_4[0:0];
  _RAND_6 = {1{`RANDOM}};
  QueueCompatibility_68_covSum = 0; //_6[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module UARTRx(
  input         clock,
  input         reset,
  input         io_en,
  input         io_in,
  output        io_out_valid,
  output [7:0]  io_out_bits,
  input  [15:0] io_div,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] debounce; // @[UARTRx.scala 24:21]
  wire  debounce_max = debounce == 2'h3; // @[UARTRx.scala 25:32]
  wire  debounce_min = debounce == 2'h0; // @[UARTRx.scala 26:32]
  reg [12:0] prescaler; // @[UARTRx.scala 28:22]
  wire  pulse = prescaler == 13'h0; // @[UARTRx.scala 30:26]
  reg [3:0] data_count; // @[UARTRx.scala 34:23]
  wire  data_last = data_count == 4'h0; // @[UARTRx.scala 35:31]
  reg [3:0] sample_count; // @[UARTRx.scala 37:25]
  wire  sample_mid = sample_count == 4'h7; // @[UARTRx.scala 38:34]
  wire [7:0] _countdown_T = {data_count,sample_count}; // @[Cat.scala 31:58]
  wire [7:0] countdown = _countdown_T - 8'h1; // @[UARTRx.scala 40:49]
  wire [3:0] remainder = io_div[3:0]; // @[UARTRx.scala 45:25]
  wire  extend = sample_count < remainder; // @[UARTRx.scala 46:30]
  reg  state; // @[UARTRx.scala 61:18]
  wire  _T_5 = ~io_in; // @[UARTRx.scala 68:13]
  wire  _GEN_8 = ~io_in & debounce_max; // @[UARTRx.scala 68:21]
  wire  start = ~state & _GEN_8; // @[UARTRx.scala 63:18]
  wire  restore = start | pulse; // @[UARTRx.scala 47:23]
  wire [12:0] prescaler_in = restore ? {{1'd0}, io_div[15:4]} : prescaler; // @[UARTRx.scala 48:25]
  wire  _prescaler_next_T_1 = restore & extend ? 1'h0 : 1'h1; // @[UARTRx.scala 49:42]
  wire [12:0] _GEN_41 = {{12'd0}, _prescaler_next_T_1}; // @[UARTRx.scala 49:37]
  wire [12:0] prescaler_next = prescaler_in - _GEN_41; // @[UARTRx.scala 49:37]
  reg [2:0] sample; // @[UARTRx.scala 51:19]
  wire  _voter_T_3 = sample[0] & sample[1]; // @[Misc.scala 166:48]
  wire  _voter_T_4 = sample[0] & sample[2]; // @[Misc.scala 166:48]
  wire  _voter_T_6 = sample[1] & sample[2]; // @[Misc.scala 166:48]
  wire  voter = _voter_T_3 | _voter_T_4 | _voter_T_6; // @[Misc.scala 167:22]
  reg [7:0] shifter; // @[UARTRx.scala 53:20]
  reg  valid; // @[UARTRx.scala 55:18]
  wire [1:0] _debounce_T_1 = debounce - 2'h1; // @[UARTRx.scala 66:30]
  wire [1:0] _GEN_0 = ~_T_5 & ~debounce_min ? _debounce_T_1 : debounce; // @[UARTRx.scala 65:41 66:18 24:21]
  wire [1:0] _debounce_T_3 = debounce + 2'h1; // @[UARTRx.scala 69:30]
  wire [3:0] _data_count_T_3 = 4'h9 - 4'h0; // @[UARTRx.scala 74:94]
  wire  _GEN_1 = debounce_max | state; // @[UARTRx.scala 70:29 71:17 61:18]
  wire [3:0] _sample_T = {sample,io_in}; // @[Cat.scala 31:58]
  wire [7:0] _shifter_T_1 = {voter,shifter[7:1]}; // @[Cat.scala 31:58]
  wire  _GEN_12 = data_last ? 1'h0 : state; // @[UARTRx.scala 102:30 103:21 61:18]
  wire [7:0] _GEN_14 = data_last ? shifter : _shifter_T_1; // @[UARTRx.scala 102:30 53:20 106:23]
  wire  _GEN_15 = sample_mid ? _GEN_12 : state; // @[UARTRx.scala 61:18 87:27]
  wire  _GEN_16 = sample_mid & data_last; // @[UARTRx.scala 87:27 56:9]
  wire [3:0] _GEN_18 = pulse ? _sample_T : {{1'd0}, sample}; // @[UARTRx.scala 82:20 83:16 51:19]
  wire  _GEN_22 = pulse & _GEN_16; // @[UARTRx.scala 82:20 56:9]
  wire [3:0] _GEN_25 = state ? _GEN_18 : {{1'd0}, sample}; // @[UARTRx.scala 63:18 51:19]
  wire [3:0] _GEN_37 = ~state ? {{1'd0}, sample} : _GEN_25; // @[UARTRx.scala 63:18 51:19]
  reg [2:0] UARTRx_covState; // @[Register tracking UARTRx state]
  reg  UARTRx_covMap [0:7]; // @[Coverage map for UARTRx]
  wire  UARTRx_covMap_read_en; // @[Coverage map for UARTRx]
  wire [2:0] UARTRx_covMap_read_addr; // @[Coverage map for UARTRx]
  wire  UARTRx_covMap_read_data; // @[Coverage map for UARTRx]
  wire  UARTRx_covMap_write_data; // @[Coverage map for UARTRx]
  wire [2:0] UARTRx_covMap_write_addr; // @[Coverage map for UARTRx]
  wire  UARTRx_covMap_write_mask; // @[Coverage map for UARTRx]
  wire  UARTRx_covMap_write_en; // @[Coverage map for UARTRx]
  reg [29:0] UARTRx_covSum; // @[Sum of coverage map]
  wire [1:0] debounce_shl;
  wire [2:0] debounce_pad;
  wire [2:0] state_shl;
  wire [2:0] state_pad;
  wire [2:0] UARTRx_xor0;
  assign io_out_valid = valid; // @[UARTRx.scala 57:16]
  assign io_out_bits = shifter; // @[UARTRx.scala 58:15]
  assign UARTRx_covMap_read_en = 1'h1;
  assign UARTRx_covMap_read_addr = UARTRx_covState;
  assign UARTRx_covMap_read_data = UARTRx_covMap[UARTRx_covMap_read_addr]; // @[Coverage map for UARTRx]
  assign UARTRx_covMap_write_data = 1'h1;
  assign UARTRx_covMap_write_addr = UARTRx_covState;
  assign UARTRx_covMap_write_mask = 1'h1;
  assign UARTRx_covMap_write_en = ~metaReset;
  assign debounce_shl = debounce;
  assign debounce_pad = {1'h0,debounce_shl};
  assign state_shl = {state, 2'h0};
  assign state_pad = state_shl;
  assign UARTRx_xor0 = debounce_pad ^ state_pad;
  assign io_covSum = UARTRx_covSum;
  always @(posedge clock) begin
    if (reset) begin // @[UARTRx.scala 24:21]
      debounce <= 2'h0; // @[UARTRx.scala 24:21]
    end else if (~io_en) begin
      debounce <= 2'h0;
    end else if (~state) begin
      if (~io_in) begin
        debounce <= _debounce_T_3;
      end else begin
        debounce <= _GEN_0;
      end
    end
    if (~state) begin // @[UARTRx.scala 63:18]
      if (~io_in) begin
        if (debounce_max) begin
          prescaler <= prescaler_next;
        end
      end
    end else if (state) begin
      prescaler <= prescaler_next;
    end
    if (~state) begin // @[UARTRx.scala 63:18]
      if (~io_in) begin
        if (debounce_max) begin
          data_count <= _data_count_T_3;
        end
      end
    end else if (state) begin
      if (pulse) begin
        data_count <= countdown[7:4];
      end
    end
    if (~state) begin // @[UARTRx.scala 63:18]
      if (~io_in) begin
        if (debounce_max) begin
          sample_count <= 4'hf;
        end
      end
    end else if (state) begin
      if (pulse) begin
        sample_count <= countdown[3:0];
      end
    end
    if (reset) begin // @[UARTRx.scala 61:18]
      state <= 1'h0; // @[UARTRx.scala 61:18]
    end else if (~state) begin
      if (~io_in) begin
        state <= _GEN_1;
      end
    end else if (state) begin
      if (pulse) begin
        state <= _GEN_15;
      end
    end
    sample <= _GEN_37[2:0];
    if (!(~state)) begin // @[UARTRx.scala 63:18]
      if (state) begin
        if (pulse) begin
          if (sample_mid) begin
            shifter <= _GEN_14;
          end
        end
      end
    end
    if (reset) begin // @[UARTRx.scala 55:18]
      valid <= 1'h0; // @[UARTRx.scala 55:18]
    end else if (~state) begin
      valid <= 1'h0;
    end else begin
      valid <= state & _GEN_22;
    end
    UARTRx_covState <= UARTRx_xor0;
    if (UARTRx_covMap_write_en & UARTRx_covMap_write_mask) begin
      UARTRx_covMap[UARTRx_covMap_write_addr] <= UARTRx_covMap_write_data; // @[Coverage map for UARTRx]
    end
    if (!(UARTRx_covMap_read_data | metaReset)) begin
      UARTRx_covSum <= UARTRx_covSum + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    UARTRx_covMap[initvar] = 0; //_9[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounce = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  prescaler = _RAND_1[12:0];
  _RAND_2 = {1{`RANDOM}};
  data_count = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  sample_count = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  sample = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  shifter = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  UARTRx_covState = 0; //_8[2:0];
  _RAND_10 = {1{`RANDOM}};
  UARTRx_covSum = 0; //_10[29:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLUART(
  input         clock,
  input         reset,
  output        auto_int_xing_out_sync_0,
  output        auto_control_xing_in_a_ready,
  input         auto_control_xing_in_a_valid,
  input  [2:0]  auto_control_xing_in_a_bits_opcode,
  input  [1:0]  auto_control_xing_in_a_bits_size,
  input  [10:0] auto_control_xing_in_a_bits_source,
  input  [30:0] auto_control_xing_in_a_bits_address,
  input  [7:0]  auto_control_xing_in_a_bits_mask,
  input  [63:0] auto_control_xing_in_a_bits_data,
  input         auto_control_xing_in_d_ready,
  output        auto_control_xing_in_d_valid,
  output [2:0]  auto_control_xing_in_d_bits_opcode,
  output [1:0]  auto_control_xing_in_d_bits_size,
  output [10:0] auto_control_xing_in_d_bits_source,
  output [63:0] auto_control_xing_in_d_bits_data,
  output        auto_io_out_txd,
  input         auto_io_out_rxd,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  buffer_auto_in_a_ready;
  wire  buffer_auto_in_a_valid;
  wire [2:0] buffer_auto_in_a_bits_opcode;
  wire [1:0] buffer_auto_in_a_bits_size;
  wire [10:0] buffer_auto_in_a_bits_source;
  wire [30:0] buffer_auto_in_a_bits_address;
  wire [7:0] buffer_auto_in_a_bits_mask;
  wire [63:0] buffer_auto_in_a_bits_data;
  wire  buffer_auto_in_d_ready;
  wire  buffer_auto_in_d_valid;
  wire [2:0] buffer_auto_in_d_bits_opcode;
  wire [1:0] buffer_auto_in_d_bits_size;
  wire [10:0] buffer_auto_in_d_bits_source;
  wire [63:0] buffer_auto_in_d_bits_data;
  wire  buffer_auto_out_a_ready;
  wire  buffer_auto_out_a_valid;
  wire [2:0] buffer_auto_out_a_bits_opcode;
  wire [1:0] buffer_auto_out_a_bits_size;
  wire [10:0] buffer_auto_out_a_bits_source;
  wire [30:0] buffer_auto_out_a_bits_address;
  wire [7:0] buffer_auto_out_a_bits_mask;
  wire [63:0] buffer_auto_out_a_bits_data;
  wire  buffer_auto_out_d_ready;
  wire  buffer_auto_out_d_valid;
  wire [2:0] buffer_auto_out_d_bits_opcode;
  wire [1:0] buffer_auto_out_d_bits_size;
  wire [10:0] buffer_auto_out_d_bits_source;
  wire [63:0] buffer_auto_out_d_bits_data;
  wire  intsource_clock; // @[Crossing.scala 26:31]
  wire  intsource_reset; // @[Crossing.scala 26:31]
  wire  intsource_auto_in_0; // @[Crossing.scala 26:31]
  wire  intsource_auto_out_sync_0; // @[Crossing.scala 26:31]
  wire [29:0] intsource_io_covSum; // @[Crossing.scala 26:31]
  wire  txm_clock; // @[UART.scala 79:19]
  wire  txm_reset; // @[UART.scala 79:19]
  wire  txm_io_en; // @[UART.scala 79:19]
  wire  txm_io_in_ready; // @[UART.scala 79:19]
  wire  txm_io_in_valid; // @[UART.scala 79:19]
  wire [7:0] txm_io_in_bits; // @[UART.scala 79:19]
  wire  txm_io_out; // @[UART.scala 79:19]
  wire [15:0] txm_io_div; // @[UART.scala 79:19]
  wire  txm_io_nstop; // @[UART.scala 79:19]
  wire [29:0] txm_io_covSum; // @[UART.scala 79:19]
  wire  txq_clock; // @[UART.scala 80:19]
  wire  txq_reset; // @[UART.scala 80:19]
  wire  txq_io_enq_ready; // @[UART.scala 80:19]
  wire  txq_io_enq_valid; // @[UART.scala 80:19]
  wire [7:0] txq_io_enq_bits; // @[UART.scala 80:19]
  wire  txq_io_deq_ready; // @[UART.scala 80:19]
  wire  txq_io_deq_valid; // @[UART.scala 80:19]
  wire [7:0] txq_io_deq_bits; // @[UART.scala 80:19]
  wire [3:0] txq_io_count; // @[UART.scala 80:19]
  wire [29:0] txq_io_covSum; // @[UART.scala 80:19]
  wire  txq_metaReset; // @[UART.scala 80:19]
  wire  rxm_clock; // @[UART.scala 82:19]
  wire  rxm_reset; // @[UART.scala 82:19]
  wire  rxm_io_en; // @[UART.scala 82:19]
  wire  rxm_io_in; // @[UART.scala 82:19]
  wire  rxm_io_out_valid; // @[UART.scala 82:19]
  wire [7:0] rxm_io_out_bits; // @[UART.scala 82:19]
  wire [15:0] rxm_io_div; // @[UART.scala 82:19]
  wire [29:0] rxm_io_covSum; // @[UART.scala 82:19]
  wire  rxm_metaReset; // @[UART.scala 82:19]
  wire  rxq_clock; // @[UART.scala 83:19]
  wire  rxq_reset; // @[UART.scala 83:19]
  wire  rxq_io_enq_ready; // @[UART.scala 83:19]
  wire  rxq_io_enq_valid; // @[UART.scala 83:19]
  wire [7:0] rxq_io_enq_bits; // @[UART.scala 83:19]
  wire  rxq_io_deq_ready; // @[UART.scala 83:19]
  wire  rxq_io_deq_valid; // @[UART.scala 83:19]
  wire [7:0] rxq_io_deq_bits; // @[UART.scala 83:19]
  wire [3:0] rxq_io_count; // @[UART.scala 83:19]
  wire [29:0] rxq_io_covSum; // @[UART.scala 83:19]
  wire  rxq_metaReset; // @[UART.scala 83:19]
  reg [15:0] div; // @[UART.scala 85:16]
  reg  txen; // @[UART.scala 91:17]
  reg  rxen; // @[UART.scala 92:17]
  reg [3:0] txwm; // @[UART.scala 99:17]
  reg [3:0] rxwm; // @[UART.scala 100:17]
  reg  nstop; // @[UART.scala 101:18]
  reg  ie_rxwm; // @[UART.scala 135:15]
  reg  ie_txwm; // @[UART.scala 135:15]
  wire  ip_txwm = txq_io_count < txwm; // @[UART.scala 138:28]
  wire  ip_rxwm = rxq_io_count > rxwm; // @[UART.scala 139:28]
  wire  _T = ~txq_io_enq_ready; // @[RegMapFIFO.scala 25:9]
  wire  _T_1 = ~rxq_io_deq_valid; // @[RegMapFIFO.scala 46:21]
  wire  in_bits_read = buffer_auto_out_a_bits_opcode == 3'h4; // @[RegisterRouter.scala 72:36]
  wire [8:0] in_bits_index = buffer_auto_out_a_bits_address[11:3]; // @[RegisterRouter.scala 71:18 73:19]
  wire [8:0] out_findex = in_bits_index & 9'h1fc; // @[RegisterRouter.scala 83:24]
  wire  _out_T = out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire [7:0] _out_backMask_T_9 = buffer_auto_out_a_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_11 = buffer_auto_out_a_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_13 = buffer_auto_out_a_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_15 = buffer_auto_out_a_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_17 = buffer_auto_out_a_bits_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_19 = buffer_auto_out_a_bits_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_21 = buffer_auto_out_a_bits_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_23 = buffer_auto_out_a_bits_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] out_backMask = {_out_backMask_T_23,_out_backMask_T_21,_out_backMask_T_19,_out_backMask_T_17,
    _out_backMask_T_15,_out_backMask_T_13,_out_backMask_T_11,_out_backMask_T_9}; // @[Cat.scala 31:58]
  wire  out_womask = &out_backMask[7:0]; // @[RegisterRouter.scala 83:24]
  wire [1:0] out_oindex = {in_bits_index[1],in_bits_index[0]}; // @[Cat.scala 31:58]
  wire [3:0] _out_backSel_T = 4'h1 << out_oindex; // @[OneHot.scala 57:35]
  wire  out_backSel_0 = _out_backSel_T[0]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_3 = buffer_auto_out_a_valid & buffer_auto_out_d_ready & in_bits_read & out_backSel_0 & out_findex
     == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_woready_0 = buffer_auto_out_a_valid & buffer_auto_out_d_ready & ~in_bits_read & out_backSel_0 & out_findex
     == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready = out_woready_0 & out_womask; // @[RegisterRouter.scala 83:24]
  wire  out_womask_2 = &out_backMask[31]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_2 = out_woready_0 & out_womask_2; // @[RegisterRouter.scala 83:24]
  wire  quash = out_f_woready_2 & buffer_auto_out_a_bits_data[31]; // @[RegMapFIFO.scala 27:26]
  wire  out_romask_3 = |out_backMask[39:32]; // @[RegisterRouter.scala 83:24]
  wire [40:0] out_prepend_3 = {1'h0,rxq_io_deq_bits,_T,31'h0}; // @[Cat.scala 31:58]
  wire [62:0] _out_T_51 = {{22'd0}, out_prepend_3}; // @[RegisterRouter.scala 83:24]
  wire [63:0] out_prepend_4 = {_T_1,_out_T_51}; // @[Cat.scala 31:58]
  wire  out_womask_6 = &out_backMask[0]; // @[RegisterRouter.scala 83:24]
  wire  out_backSel_1 = _out_backSel_T[1]; // @[RegisterRouter.scala 83:24]
  wire  out_woready_6 = buffer_auto_out_a_valid & buffer_auto_out_d_ready & ~in_bits_read & out_backSel_1 & out_findex
     == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_6 = out_woready_6 & out_womask_6; // @[RegisterRouter.scala 83:24]
  wire  out_womask_7 = &out_backMask[1]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_7 = out_woready_6 & out_womask_7; // @[RegisterRouter.scala 83:24]
  wire [1:0] out_prepend_5 = {nstop,txen}; // @[Cat.scala 31:58]
  wire  out_womask_8 = &out_backMask[19:16]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_8 = out_woready_6 & out_womask_8; // @[RegisterRouter.scala 83:24]
  wire [15:0] _out_prepend_T_6 = {{14'd0}, out_prepend_5}; // @[RegisterRouter.scala 83:24]
  wire [19:0] out_prepend_6 = {txwm,_out_prepend_T_6}; // @[Cat.scala 31:58]
  wire  out_womask_9 = &out_backMask[32]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_9 = out_woready_6 & out_womask_9; // @[RegisterRouter.scala 83:24]
  wire [31:0] _out_prepend_T_7 = {{12'd0}, out_prepend_6}; // @[RegisterRouter.scala 83:24]
  wire [32:0] out_prepend_7 = {rxen,_out_prepend_T_7}; // @[Cat.scala 31:58]
  wire  out_womask_10 = &out_backMask[51:48]; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_10 = out_woready_6 & out_womask_10; // @[RegisterRouter.scala 83:24]
  wire [47:0] _out_prepend_T_8 = {{15'd0}, out_prepend_7}; // @[RegisterRouter.scala 83:24]
  wire [51:0] out_prepend_8 = {rxwm,_out_prepend_T_8}; // @[Cat.scala 31:58]
  wire  out_backSel_2 = _out_backSel_T[2]; // @[RegisterRouter.scala 83:24]
  wire  out_woready_11 = buffer_auto_out_a_valid & buffer_auto_out_d_ready & ~in_bits_read & out_backSel_2 & out_findex
     == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_11 = out_woready_11 & out_womask_6; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_12 = out_woready_11 & out_womask_7; // @[RegisterRouter.scala 83:24]
  wire [1:0] out_prepend_9 = {ie_rxwm,ie_txwm}; // @[Cat.scala 31:58]
  wire [31:0] _out_prepend_T_10 = {{30'd0}, out_prepend_9}; // @[RegisterRouter.scala 83:24]
  wire [33:0] out_prepend_11 = {ip_rxwm,ip_txwm,_out_prepend_T_10}; // @[Cat.scala 31:58]
  wire  out_womask_15 = &out_backMask[15:0]; // @[RegisterRouter.scala 83:24]
  wire  out_backSel_3 = _out_backSel_T[3]; // @[RegisterRouter.scala 83:24]
  wire  out_woready_15 = buffer_auto_out_a_valid & buffer_auto_out_d_ready & ~in_bits_read & out_backSel_3 & out_findex
     == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_woready_15 = out_woready_15 & out_womask_15; // @[RegisterRouter.scala 83:24]
  wire  _GEN_25 = 2'h1 == out_oindex ? _out_T : _out_T; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_26 = 2'h2 == out_oindex ? _out_T : _GEN_25; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_27 = 2'h3 == out_oindex ? _out_T : _GEN_26; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _out_out_bits_data_WIRE_1_1 = {{12'd0}, out_prepend_8}; // @[MuxLiteral.scala 48:{48,48}]
  wire [63:0] _GEN_29 = 2'h1 == out_oindex ? _out_out_bits_data_WIRE_1_1 : out_prepend_4; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _out_out_bits_data_WIRE_1_2 = {{30'd0}, out_prepend_11}; // @[MuxLiteral.scala 48:{48,48}]
  wire [63:0] _GEN_30 = 2'h2 == out_oindex ? _out_out_bits_data_WIRE_1_2 : _GEN_29; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _out_out_bits_data_WIRE_1_3 = {{48'd0}, div}; // @[MuxLiteral.scala 48:{48,48}]
  wire [63:0] _GEN_31 = 2'h3 == out_oindex ? _out_out_bits_data_WIRE_1_3 : _GEN_30; // @[MuxLiteral.scala 48:{10,10}]
  wire [29:0] TLUART_covSum;
  wire [29:0] txq_sum;
  wire [29:0] rxq_sum;
  wire [29:0] txm_sum;
  wire [29:0] intsource_sum;
  wire [29:0] rxm_sum;
  IntSyncCrossingSource_1 intsource ( // @[Crossing.scala 26:31]
    .clock(intsource_clock),
    .reset(intsource_reset),
    .auto_in_0(intsource_auto_in_0),
    .auto_out_sync_0(intsource_auto_out_sync_0),
    .io_covSum(intsource_io_covSum)
  );
  UARTTx txm ( // @[UART.scala 79:19]
    .clock(txm_clock),
    .reset(txm_reset),
    .io_en(txm_io_en),
    .io_in_ready(txm_io_in_ready),
    .io_in_valid(txm_io_in_valid),
    .io_in_bits(txm_io_in_bits),
    .io_out(txm_io_out),
    .io_div(txm_io_div),
    .io_nstop(txm_io_nstop),
    .io_covSum(txm_io_covSum)
  );
  QueueCompatibility_68 txq ( // @[UART.scala 80:19]
    .clock(txq_clock),
    .reset(txq_reset),
    .io_enq_ready(txq_io_enq_ready),
    .io_enq_valid(txq_io_enq_valid),
    .io_enq_bits(txq_io_enq_bits),
    .io_deq_ready(txq_io_deq_ready),
    .io_deq_valid(txq_io_deq_valid),
    .io_deq_bits(txq_io_deq_bits),
    .io_count(txq_io_count),
    .io_covSum(txq_io_covSum),
    .metaReset(txq_metaReset)
  );
  UARTRx rxm ( // @[UART.scala 82:19]
    .clock(rxm_clock),
    .reset(rxm_reset),
    .io_en(rxm_io_en),
    .io_in(rxm_io_in),
    .io_out_valid(rxm_io_out_valid),
    .io_out_bits(rxm_io_out_bits),
    .io_div(rxm_io_div),
    .io_covSum(rxm_io_covSum),
    .metaReset(rxm_metaReset)
  );
  QueueCompatibility_68 rxq ( // @[UART.scala 83:19]
    .clock(rxq_clock),
    .reset(rxq_reset),
    .io_enq_ready(rxq_io_enq_ready),
    .io_enq_valid(rxq_io_enq_valid),
    .io_enq_bits(rxq_io_enq_bits),
    .io_deq_ready(rxq_io_deq_ready),
    .io_deq_valid(rxq_io_deq_valid),
    .io_deq_bits(rxq_io_deq_bits),
    .io_count(rxq_io_count),
    .io_covSum(rxq_io_covSum),
    .metaReset(rxq_metaReset)
  );
  assign buffer_auto_in_a_ready = buffer_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_valid = buffer_auto_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_opcode = buffer_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_size = buffer_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_source = buffer_auto_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_in_d_bits_data = buffer_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign buffer_auto_out_a_valid = buffer_auto_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_opcode = buffer_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_size = buffer_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_source = buffer_auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_address = buffer_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_mask = buffer_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_bits_data = buffer_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_d_ready = buffer_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_int_xing_out_sync_0 = intsource_auto_out_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_control_xing_in_a_ready = buffer_auto_in_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_control_xing_in_d_valid = buffer_auto_in_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_control_xing_in_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_control_xing_in_d_bits_size = buffer_auto_in_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_control_xing_in_d_bits_source = buffer_auto_in_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_control_xing_in_d_bits_data = buffer_auto_in_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign auto_io_out_txd = txm_io_out; // @[Nodes.scala 1207:84 UART.scala 113:12]
  assign buffer_auto_in_a_valid = auto_control_xing_in_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_opcode = auto_control_xing_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_size = auto_control_xing_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_source = auto_control_xing_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_address = auto_control_xing_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_mask = auto_control_xing_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_a_bits_data = auto_control_xing_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_in_d_ready = auto_control_xing_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign buffer_auto_out_a_ready = buffer_auto_out_d_ready; // @[RegisterRouter.scala 83:24]
  assign buffer_auto_out_d_valid = buffer_auto_out_a_valid; // @[RegisterRouter.scala 83:24]
  assign buffer_auto_out_d_bits_opcode = {{2'd0}, in_bits_read}; // @[Nodes.scala 1210:84 RegisterRouter.scala 98:19]
  assign buffer_auto_out_d_bits_size = buffer_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_source = buffer_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign buffer_auto_out_d_bits_data = _GEN_27 ? _GEN_31 : 64'h0; // @[RegisterRouter.scala 83:24]
  assign intsource_clock = clock;
  assign intsource_reset = reset;
  assign intsource_auto_in_0 = ip_txwm & ie_txwm | ip_rxwm & ie_rxwm; // @[UART.scala 140:41]
  assign txm_clock = clock;
  assign txm_reset = reset;
  assign txm_io_en = txen; // @[UART.scala 109:15]
  assign txm_io_in_valid = txq_io_deq_valid; // @[UART.scala 110:13]
  assign txm_io_in_bits = txq_io_deq_bits; // @[UART.scala 110:13]
  assign txm_io_div = div; // @[UART.scala 111:14]
  assign txm_io_nstop = nstop; // @[UART.scala 112:16]
  assign txq_clock = clock;
  assign txq_reset = reset;
  assign txq_io_enq_valid = out_f_woready & ~quash; // @[RegMapFIFO.scala 19:30]
  assign txq_io_enq_bits = buffer_auto_out_a_bits_data[7:0]; // @[RegisterRouter.scala 83:24]
  assign txq_io_deq_ready = txm_io_in_ready; // @[UART.scala 110:13]
  assign rxm_clock = clock;
  assign rxm_reset = reset;
  assign rxm_io_en = rxen; // @[UART.scala 120:13]
  assign rxm_io_in = auto_io_out_rxd; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign rxm_io_div = div; // @[UART.scala 123:14]
  assign rxq_clock = clock;
  assign rxq_reset = reset;
  assign rxq_io_enq_valid = rxm_io_out_valid; // @[UART.scala 122:14]
  assign rxq_io_enq_bits = rxm_io_out_bits; // @[UART.scala 122:14]
  assign rxq_io_deq_ready = out_roready_3 & out_romask_3; // @[RegisterRouter.scala 83:24]
  assign TLUART_covSum = 30'h0;
  assign txq_sum = TLUART_covSum + txq_io_covSum;
  assign rxq_sum = txq_sum + rxq_io_covSum;
  assign txm_sum = rxq_sum + txm_io_covSum;
  assign intsource_sum = txm_sum + intsource_io_covSum;
  assign rxm_sum = intsource_sum + rxm_io_covSum;
  assign io_covSum = rxm_sum;
  assign txq_metaReset = metaReset;
  assign rxq_metaReset = metaReset;
  assign rxm_metaReset = metaReset;
  always @(posedge clock) begin
    if (reset) begin // @[UART.scala 85:16]
      div <= 16'h364; // @[UART.scala 85:16]
    end else if (out_f_woready_15) begin
      div <= buffer_auto_out_a_bits_data[15:0];
    end
    if (reset) begin // @[UART.scala 91:17]
      txen <= 1'h0; // @[UART.scala 91:17]
    end else if (out_f_woready_6) begin
      txen <= buffer_auto_out_a_bits_data[0];
    end
    if (reset) begin // @[UART.scala 92:17]
      rxen <= 1'h0; // @[UART.scala 92:17]
    end else if (out_f_woready_9) begin
      rxen <= buffer_auto_out_a_bits_data[32];
    end
    if (reset) begin // @[UART.scala 99:17]
      txwm <= 4'h0; // @[UART.scala 99:17]
    end else if (out_f_woready_8) begin
      txwm <= buffer_auto_out_a_bits_data[19:16];
    end
    if (reset) begin // @[UART.scala 100:17]
      rxwm <= 4'h0; // @[UART.scala 100:17]
    end else if (out_f_woready_10) begin
      rxwm <= buffer_auto_out_a_bits_data[51:48];
    end
    if (reset) begin // @[UART.scala 101:18]
      nstop <= 1'h0; // @[UART.scala 101:18]
    end else if (out_f_woready_7) begin
      nstop <= buffer_auto_out_a_bits_data[1];
    end
    if (reset) begin // @[UART.scala 135:15]
      ie_rxwm <= 1'h0; // @[UART.scala 135:15]
    end else if (out_f_woready_12) begin
      ie_rxwm <= buffer_auto_out_a_bits_data[1];
    end
    if (reset) begin // @[UART.scala 135:15]
      ie_txwm <= 1'h0; // @[UART.scala 135:15]
    end else if (out_f_woready_11) begin
      ie_txwm <= buffer_auto_out_a_bits_data[0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  div = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  txen = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  rxen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  txwm = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  rxwm = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  nstop = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  ie_rxwm = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  ie_txwm = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain_2(
  output        auto_uart_0_int_xing_out_sync_0,
  output        auto_uart_0_control_xing_in_a_ready,
  input         auto_uart_0_control_xing_in_a_valid,
  input  [2:0]  auto_uart_0_control_xing_in_a_bits_opcode,
  input  [1:0]  auto_uart_0_control_xing_in_a_bits_size,
  input  [10:0] auto_uart_0_control_xing_in_a_bits_source,
  input  [30:0] auto_uart_0_control_xing_in_a_bits_address,
  input  [7:0]  auto_uart_0_control_xing_in_a_bits_mask,
  input  [63:0] auto_uart_0_control_xing_in_a_bits_data,
  input         auto_uart_0_control_xing_in_d_ready,
  output        auto_uart_0_control_xing_in_d_valid,
  output [2:0]  auto_uart_0_control_xing_in_d_bits_opcode,
  output [1:0]  auto_uart_0_control_xing_in_d_bits_size,
  output [10:0] auto_uart_0_control_xing_in_d_bits_source,
  output [63:0] auto_uart_0_control_xing_in_d_bits_data,
  output        auto_uart_0_io_out_txd,
  input         auto_uart_0_io_out_rxd,
  input         auto_clock_in_clock,
  input         auto_clock_in_reset,
  output [29:0] io_covSum,
  input         metaReset
);
  wire  uart_0_clock; // @[UART.scala 243:51]
  wire  uart_0_reset; // @[UART.scala 243:51]
  wire  uart_0_auto_int_xing_out_sync_0; // @[UART.scala 243:51]
  wire  uart_0_auto_control_xing_in_a_ready; // @[UART.scala 243:51]
  wire  uart_0_auto_control_xing_in_a_valid; // @[UART.scala 243:51]
  wire [2:0] uart_0_auto_control_xing_in_a_bits_opcode; // @[UART.scala 243:51]
  wire [1:0] uart_0_auto_control_xing_in_a_bits_size; // @[UART.scala 243:51]
  wire [10:0] uart_0_auto_control_xing_in_a_bits_source; // @[UART.scala 243:51]
  wire [30:0] uart_0_auto_control_xing_in_a_bits_address; // @[UART.scala 243:51]
  wire [7:0] uart_0_auto_control_xing_in_a_bits_mask; // @[UART.scala 243:51]
  wire [63:0] uart_0_auto_control_xing_in_a_bits_data; // @[UART.scala 243:51]
  wire  uart_0_auto_control_xing_in_d_ready; // @[UART.scala 243:51]
  wire  uart_0_auto_control_xing_in_d_valid; // @[UART.scala 243:51]
  wire [2:0] uart_0_auto_control_xing_in_d_bits_opcode; // @[UART.scala 243:51]
  wire [1:0] uart_0_auto_control_xing_in_d_bits_size; // @[UART.scala 243:51]
  wire [10:0] uart_0_auto_control_xing_in_d_bits_source; // @[UART.scala 243:51]
  wire [63:0] uart_0_auto_control_xing_in_d_bits_data; // @[UART.scala 243:51]
  wire  uart_0_auto_io_out_txd; // @[UART.scala 243:51]
  wire  uart_0_auto_io_out_rxd; // @[UART.scala 243:51]
  wire [29:0] uart_0_io_covSum; // @[UART.scala 243:51]
  wire  uart_0_metaReset; // @[UART.scala 243:51]
  wire [29:0] ClockSinkDomain_2_covSum;
  wire [29:0] uart_0_sum;
  TLUART uart_0 ( // @[UART.scala 243:51]
    .clock(uart_0_clock),
    .reset(uart_0_reset),
    .auto_int_xing_out_sync_0(uart_0_auto_int_xing_out_sync_0),
    .auto_control_xing_in_a_ready(uart_0_auto_control_xing_in_a_ready),
    .auto_control_xing_in_a_valid(uart_0_auto_control_xing_in_a_valid),
    .auto_control_xing_in_a_bits_opcode(uart_0_auto_control_xing_in_a_bits_opcode),
    .auto_control_xing_in_a_bits_size(uart_0_auto_control_xing_in_a_bits_size),
    .auto_control_xing_in_a_bits_source(uart_0_auto_control_xing_in_a_bits_source),
    .auto_control_xing_in_a_bits_address(uart_0_auto_control_xing_in_a_bits_address),
    .auto_control_xing_in_a_bits_mask(uart_0_auto_control_xing_in_a_bits_mask),
    .auto_control_xing_in_a_bits_data(uart_0_auto_control_xing_in_a_bits_data),
    .auto_control_xing_in_d_ready(uart_0_auto_control_xing_in_d_ready),
    .auto_control_xing_in_d_valid(uart_0_auto_control_xing_in_d_valid),
    .auto_control_xing_in_d_bits_opcode(uart_0_auto_control_xing_in_d_bits_opcode),
    .auto_control_xing_in_d_bits_size(uart_0_auto_control_xing_in_d_bits_size),
    .auto_control_xing_in_d_bits_source(uart_0_auto_control_xing_in_d_bits_source),
    .auto_control_xing_in_d_bits_data(uart_0_auto_control_xing_in_d_bits_data),
    .auto_io_out_txd(uart_0_auto_io_out_txd),
    .auto_io_out_rxd(uart_0_auto_io_out_rxd),
    .io_covSum(uart_0_io_covSum),
    .metaReset(uart_0_metaReset)
  );
  assign auto_uart_0_int_xing_out_sync_0 = uart_0_auto_int_xing_out_sync_0; // @[LazyModule.scala 311:12]
  assign auto_uart_0_control_xing_in_a_ready = uart_0_auto_control_xing_in_a_ready; // @[LazyModule.scala 309:16]
  assign auto_uart_0_control_xing_in_d_valid = uart_0_auto_control_xing_in_d_valid; // @[LazyModule.scala 309:16]
  assign auto_uart_0_control_xing_in_d_bits_opcode = uart_0_auto_control_xing_in_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign auto_uart_0_control_xing_in_d_bits_size = uart_0_auto_control_xing_in_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_uart_0_control_xing_in_d_bits_source = uart_0_auto_control_xing_in_d_bits_source; // @[LazyModule.scala 309:16]
  assign auto_uart_0_control_xing_in_d_bits_data = uart_0_auto_control_xing_in_d_bits_data; // @[LazyModule.scala 309:16]
  assign auto_uart_0_io_out_txd = uart_0_auto_io_out_txd; // @[LazyModule.scala 311:12]
  assign uart_0_clock = auto_clock_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign uart_0_reset = auto_clock_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign uart_0_auto_control_xing_in_a_valid = auto_uart_0_control_xing_in_a_valid; // @[LazyModule.scala 309:16]
  assign uart_0_auto_control_xing_in_a_bits_opcode = auto_uart_0_control_xing_in_a_bits_opcode; // @[LazyModule.scala 309:16]
  assign uart_0_auto_control_xing_in_a_bits_size = auto_uart_0_control_xing_in_a_bits_size; // @[LazyModule.scala 309:16]
  assign uart_0_auto_control_xing_in_a_bits_source = auto_uart_0_control_xing_in_a_bits_source; // @[LazyModule.scala 309:16]
  assign uart_0_auto_control_xing_in_a_bits_address = auto_uart_0_control_xing_in_a_bits_address; // @[LazyModule.scala 309:16]
  assign uart_0_auto_control_xing_in_a_bits_mask = auto_uart_0_control_xing_in_a_bits_mask; // @[LazyModule.scala 309:16]
  assign uart_0_auto_control_xing_in_a_bits_data = auto_uart_0_control_xing_in_a_bits_data; // @[LazyModule.scala 309:16]
  assign uart_0_auto_control_xing_in_d_ready = auto_uart_0_control_xing_in_d_ready; // @[LazyModule.scala 309:16]
  assign uart_0_auto_io_out_rxd = auto_uart_0_io_out_rxd; // @[LazyModule.scala 311:12]
  assign ClockSinkDomain_2_covSum = 30'h0;
  assign uart_0_sum = ClockSinkDomain_2_covSum + uart_0_io_covSum;
  assign io_covSum = uart_0_sum;
  assign uart_0_metaReset = metaReset;
endmodule
module MagicDevice(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [1:0]  auto_in_a_bits_size,
  input  [10:0] auto_in_a_bits_source,
  input  [11:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_size,
  output [10:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  output [29:0] io_covSum
);
  wire  impl_clock; // @[Magic.scala 69:22]
  wire  impl_reset; // @[Magic.scala 69:22]
  wire [11:0] impl_read_select; // @[Magic.scala 69:22]
  wire  impl_read_ready; // @[Magic.scala 69:22]
  wire  impl_read_valid; // @[Magic.scala 69:22]
  wire [63:0] impl_read_data; // @[Magic.scala 69:22]
  wire  in_bits_read = auto_in_a_bits_opcode == 3'h4; // @[RegisterRouter.scala 72:36]
  wire [8:0] in_bits_index = auto_in_a_bits_address[11:3]; // @[Edges.scala 191:34]
  wire [3:0] out_iindex = {in_bits_index[3],in_bits_index[2],in_bits_index[1],in_bits_index[0]}; // @[Cat.scala 31:58]
  wire [8:0] out_findex = in_bits_index & 9'h1f0; // @[RegisterRouter.scala 83:24]
  wire  _out_T_14 = out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire [15:0] _out_backSel_T = 16'h1 << out_iindex; // @[OneHot.scala 57:35]
  wire  out_backSel_0 = _out_backSel_T[0]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_0 = auto_in_a_valid & auto_in_d_ready & in_bits_read & out_backSel_0 & out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire [7:0] _out_backMask_T_23 = auto_in_a_bits_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_21 = auto_in_a_bits_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_19 = auto_in_a_bits_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_17 = auto_in_a_bits_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_15 = auto_in_a_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_13 = auto_in_a_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_11 = auto_in_a_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_9 = auto_in_a_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] out_backMask = {_out_backMask_T_23,_out_backMask_T_21,_out_backMask_T_19,_out_backMask_T_17,
    _out_backMask_T_15,_out_backMask_T_13,_out_backMask_T_11,_out_backMask_T_9}; // @[Cat.scala 31:58]
  wire  out_romask = |out_backMask; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready = out_roready_0 & out_romask; // @[RegisterRouter.scala 83:24]
  wire  out_backSel_1 = _out_backSel_T[1]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_2 = auto_in_a_valid & auto_in_d_ready & in_bits_read & out_backSel_1 & out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_2 = out_roready_2 & out_romask; // @[RegisterRouter.scala 83:24]
  wire [11:0] _GEN_1 = out_f_roready_2 ? 12'h8 : 12'h0; // @[Magic.scala 76:22 77:29]
  wire  out_backSel_2 = _out_backSel_T[2]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_4 = auto_in_a_valid & auto_in_d_ready & in_bits_read & out_backSel_2 & out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_4 = out_roready_4 & out_romask; // @[RegisterRouter.scala 83:24]
  wire [11:0] _GEN_2 = out_f_roready_4 ? 12'h10 : _GEN_1; // @[Magic.scala 76:22 77:29]
  wire  out_backSel_3 = _out_backSel_T[3]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_6 = auto_in_a_valid & auto_in_d_ready & in_bits_read & out_backSel_3 & out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_6 = out_roready_6 & out_romask; // @[RegisterRouter.scala 83:24]
  wire [11:0] _GEN_3 = out_f_roready_6 ? 12'h18 : _GEN_2; // @[Magic.scala 76:22 77:29]
  wire  out_backSel_4 = _out_backSel_T[4]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_8 = auto_in_a_valid & auto_in_d_ready & in_bits_read & out_backSel_4 & out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_8 = out_roready_8 & out_romask; // @[RegisterRouter.scala 83:24]
  wire [11:0] _GEN_4 = out_f_roready_8 ? 12'h20 : _GEN_3; // @[Magic.scala 76:22 77:29]
  wire  out_backSel_5 = _out_backSel_T[5]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_1 = auto_in_a_valid & auto_in_d_ready & in_bits_read & out_backSel_5 & out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_1 = out_roready_1 & out_romask; // @[RegisterRouter.scala 83:24]
  wire [11:0] _GEN_5 = out_f_roready_1 ? 12'h28 : _GEN_4; // @[Magic.scala 76:22 77:29]
  wire  out_backSel_6 = _out_backSel_T[6]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_3 = auto_in_a_valid & auto_in_d_ready & in_bits_read & out_backSel_6 & out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_3 = out_roready_3 & out_romask; // @[RegisterRouter.scala 83:24]
  wire [11:0] _GEN_6 = out_f_roready_3 ? 12'h30 : _GEN_5; // @[Magic.scala 76:22 77:29]
  wire  out_backSel_7 = _out_backSel_T[7]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_5 = auto_in_a_valid & auto_in_d_ready & in_bits_read & out_backSel_7 & out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_5 = out_roready_5 & out_romask; // @[RegisterRouter.scala 83:24]
  wire [11:0] _GEN_7 = out_f_roready_5 ? 12'h38 : _GEN_6; // @[Magic.scala 76:22 77:29]
  wire  out_backSel_8 = _out_backSel_T[8]; // @[RegisterRouter.scala 83:24]
  wire  out_roready_7 = auto_in_a_valid & auto_in_d_ready & in_bits_read & out_backSel_8 & out_findex == 9'h0; // @[RegisterRouter.scala 83:24]
  wire  out_f_roready_7 = out_roready_7 & out_romask; // @[RegisterRouter.scala 83:24]
  wire  field_wire_8_valid = impl_read_valid; // @[Magic.scala 64:48 75:16]
  wire  out_rofireMux_out_8 = field_wire_8_valid | ~out_romask; // @[RegisterRouter.scala 83:24]
  wire  _out_rofireMux_T_37 = out_rofireMux_out_8 | ~(out_findex == 9'h0); // @[RegisterRouter.scala 83:24]
  wire  _GEN_42 = 4'h1 == out_iindex ? _out_rofireMux_T_37 : _out_rofireMux_T_37; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_43 = 4'h2 == out_iindex ? _out_rofireMux_T_37 : _GEN_42; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_44 = 4'h3 == out_iindex ? _out_rofireMux_T_37 : _GEN_43; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_45 = 4'h4 == out_iindex ? _out_rofireMux_T_37 : _GEN_44; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_46 = 4'h5 == out_iindex ? _out_rofireMux_T_37 : _GEN_45; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_47 = 4'h6 == out_iindex ? _out_rofireMux_T_37 : _GEN_46; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_48 = 4'h7 == out_iindex ? _out_rofireMux_T_37 : _GEN_47; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_49 = 4'h8 == out_iindex ? _out_rofireMux_T_37 : _GEN_48; // @[MuxLiteral.scala 48:{10,10}]
  wire  out_rofireMux = 4'hf == out_iindex | (4'he == out_iindex | (4'hd == out_iindex | (4'hc == out_iindex | (4'hb ==
    out_iindex | (4'ha == out_iindex | (4'h9 == out_iindex | _GEN_49)))))); // @[MuxLiteral.scala 48:{10,10}]
  wire  out_oready = in_bits_read ? out_rofireMux : 1'h1; // @[RegisterRouter.scala 83:24]
  wire [63:0] field_wire_0_bits = impl_read_data; // @[Magic.scala 64:48 74:15]
  wire  _GEN_74 = 4'h1 == out_iindex ? _out_T_14 : _out_T_14; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_75 = 4'h2 == out_iindex ? _out_T_14 : _GEN_74; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_76 = 4'h3 == out_iindex ? _out_T_14 : _GEN_75; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_77 = 4'h4 == out_iindex ? _out_T_14 : _GEN_76; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_78 = 4'h5 == out_iindex ? _out_T_14 : _GEN_77; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_79 = 4'h6 == out_iindex ? _out_T_14 : _GEN_78; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_80 = 4'h7 == out_iindex ? _out_T_14 : _GEN_79; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_81 = 4'h8 == out_iindex ? _out_T_14 : _GEN_80; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_88 = 4'hf == out_iindex | (4'he == out_iindex | (4'hd == out_iindex | (4'hc == out_iindex | (4'hb ==
    out_iindex | (4'ha == out_iindex | (4'h9 == out_iindex | _GEN_81)))))); // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_90 = 4'h1 == out_iindex ? field_wire_0_bits : field_wire_0_bits; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_91 = 4'h2 == out_iindex ? field_wire_0_bits : _GEN_90; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_92 = 4'h3 == out_iindex ? field_wire_0_bits : _GEN_91; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_93 = 4'h4 == out_iindex ? field_wire_0_bits : _GEN_92; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_94 = 4'h5 == out_iindex ? field_wire_0_bits : _GEN_93; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_95 = 4'h6 == out_iindex ? field_wire_0_bits : _GEN_94; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_96 = 4'h7 == out_iindex ? field_wire_0_bits : _GEN_95; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_97 = 4'h8 == out_iindex ? field_wire_0_bits : _GEN_96; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_98 = 4'h9 == out_iindex ? 64'h0 : _GEN_97; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_99 = 4'ha == out_iindex ? 64'h0 : _GEN_98; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_100 = 4'hb == out_iindex ? 64'h0 : _GEN_99; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_101 = 4'hc == out_iindex ? 64'h0 : _GEN_100; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_102 = 4'hd == out_iindex ? 64'h0 : _GEN_101; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_103 = 4'he == out_iindex ? 64'h0 : _GEN_102; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_104 = 4'hf == out_iindex ? 64'h0 : _GEN_103; // @[MuxLiteral.scala 48:{10,10}]
  wire [29:0] MagicDevice_covSum;
  MagicDeviceBlackbox impl ( // @[Magic.scala 69:22]
    .clock(impl_clock),
    .reset(impl_reset),
    .read_select(impl_read_select),
    .read_ready(impl_read_ready),
    .read_valid(impl_read_valid),
    .read_data(impl_read_data)
  );
  assign auto_in_a_ready = auto_in_d_ready & out_oready; // @[RegisterRouter.scala 83:24]
  assign auto_in_d_valid = auto_in_a_valid & out_oready; // @[RegisterRouter.scala 83:24]
  assign auto_in_d_bits_opcode = {{2'd0}, in_bits_read}; // @[Nodes.scala 1210:84 RegisterRouter.scala 98:19]
  assign auto_in_d_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_in_d_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_in_d_bits_data = _GEN_88 ? _GEN_104 : 64'h0; // @[RegisterRouter.scala 83:24]
  assign impl_clock = clock; // @[Magic.scala 70:19]
  assign impl_reset = reset; // @[Magic.scala 71:28]
  assign impl_read_select = out_f_roready_7 ? 12'h40 : _GEN_7; // @[Magic.scala 76:22 77:29]
  assign impl_read_ready = out_f_roready | out_f_roready_2 | out_f_roready_4 | out_f_roready_6 | out_f_roready_8 |
    out_f_roready_1 | out_f_roready_3 | out_f_roready_5 | out_f_roready_7; // @[Magic.scala 81:73]
  assign MagicDevice_covSum = 30'h0;
  assign io_covSum = MagicDevice_covSum;
endmodule
module StarshipASICTop(
  input         clock,
  input         reset,
  input         mem_axi4_0_aw_ready,
  output        mem_axi4_0_aw_valid,
  output [3:0]  mem_axi4_0_aw_bits_id,
  output [31:0] mem_axi4_0_aw_bits_addr,
  output [7:0]  mem_axi4_0_aw_bits_len,
  output [2:0]  mem_axi4_0_aw_bits_size,
  output [1:0]  mem_axi4_0_aw_bits_burst,
  output        mem_axi4_0_aw_bits_lock,
  output [3:0]  mem_axi4_0_aw_bits_cache,
  output [2:0]  mem_axi4_0_aw_bits_prot,
  output [3:0]  mem_axi4_0_aw_bits_qos,
  input         mem_axi4_0_w_ready,
  output        mem_axi4_0_w_valid,
  output [63:0] mem_axi4_0_w_bits_data,
  output [7:0]  mem_axi4_0_w_bits_strb,
  output        mem_axi4_0_w_bits_last,
  output        mem_axi4_0_b_ready,
  input         mem_axi4_0_b_valid,
  input  [3:0]  mem_axi4_0_b_bits_id,
  input  [1:0]  mem_axi4_0_b_bits_resp,
  input         mem_axi4_0_ar_ready,
  output        mem_axi4_0_ar_valid,
  output [3:0]  mem_axi4_0_ar_bits_id,
  output [31:0] mem_axi4_0_ar_bits_addr,
  output [7:0]  mem_axi4_0_ar_bits_len,
  output [2:0]  mem_axi4_0_ar_bits_size,
  output [1:0]  mem_axi4_0_ar_bits_burst,
  output        mem_axi4_0_ar_bits_lock,
  output [3:0]  mem_axi4_0_ar_bits_cache,
  output [2:0]  mem_axi4_0_ar_bits_prot,
  output [3:0]  mem_axi4_0_ar_bits_qos,
  output        mem_axi4_0_r_ready,
  input         mem_axi4_0_r_valid,
  input  [3:0]  mem_axi4_0_r_bits_id,
  input  [63:0] mem_axi4_0_r_bits_data,
  input  [1:0]  mem_axi4_0_r_bits_resp,
  input         mem_axi4_0_r_bits_last,
  output        l2_frontend_bus_axi4_0_aw_ready,
  input         l2_frontend_bus_axi4_0_aw_valid,
  input  [7:0]  l2_frontend_bus_axi4_0_aw_bits_id,
  input  [31:0] l2_frontend_bus_axi4_0_aw_bits_addr,
  input  [7:0]  l2_frontend_bus_axi4_0_aw_bits_len,
  input  [2:0]  l2_frontend_bus_axi4_0_aw_bits_size,
  input  [1:0]  l2_frontend_bus_axi4_0_aw_bits_burst,
  input         l2_frontend_bus_axi4_0_aw_bits_lock,
  input  [3:0]  l2_frontend_bus_axi4_0_aw_bits_cache,
  input  [2:0]  l2_frontend_bus_axi4_0_aw_bits_prot,
  input  [3:0]  l2_frontend_bus_axi4_0_aw_bits_qos,
  output        l2_frontend_bus_axi4_0_w_ready,
  input         l2_frontend_bus_axi4_0_w_valid,
  input  [63:0] l2_frontend_bus_axi4_0_w_bits_data,
  input  [7:0]  l2_frontend_bus_axi4_0_w_bits_strb,
  input         l2_frontend_bus_axi4_0_w_bits_last,
  input         l2_frontend_bus_axi4_0_b_ready,
  output        l2_frontend_bus_axi4_0_b_valid,
  output [7:0]  l2_frontend_bus_axi4_0_b_bits_id,
  output [1:0]  l2_frontend_bus_axi4_0_b_bits_resp,
  output        l2_frontend_bus_axi4_0_ar_ready,
  input         l2_frontend_bus_axi4_0_ar_valid,
  input  [7:0]  l2_frontend_bus_axi4_0_ar_bits_id,
  input  [31:0] l2_frontend_bus_axi4_0_ar_bits_addr,
  input  [7:0]  l2_frontend_bus_axi4_0_ar_bits_len,
  input  [2:0]  l2_frontend_bus_axi4_0_ar_bits_size,
  input  [1:0]  l2_frontend_bus_axi4_0_ar_bits_burst,
  input         l2_frontend_bus_axi4_0_ar_bits_lock,
  input  [3:0]  l2_frontend_bus_axi4_0_ar_bits_cache,
  input  [2:0]  l2_frontend_bus_axi4_0_ar_bits_prot,
  input  [3:0]  l2_frontend_bus_axi4_0_ar_bits_qos,
  input         l2_frontend_bus_axi4_0_r_ready,
  output        l2_frontend_bus_axi4_0_r_valid,
  output [7:0]  l2_frontend_bus_axi4_0_r_bits_id,
  output [63:0] l2_frontend_bus_axi4_0_r_bits_data,
  output [1:0]  l2_frontend_bus_axi4_0_r_bits_resp,
  output        l2_frontend_bus_axi4_0_r_bits_last,
  output        uart_0_txd,
  input         uart_0_rxd,
  output [29:0] io_covSum,
  input         metaReset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  ibus_auto_int_bus_int_in_0;
  wire  ibus_auto_int_bus_int_out_0;
  wire  ibus_int_bus_auto_int_in_0; // @[InterruptBus.scala 14:27]
  wire  ibus_int_bus_auto_int_out_0; // @[InterruptBus.scala 14:27]
  wire [29:0] ibus_int_bus_io_covSum; // @[InterruptBus.scala 14:27]
  wire  dummyClockGroupSourceNode_clock; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_reset; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_clock; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_reset; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_clock; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_reset; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_clock; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_reset; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_clock; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_reset; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_clock; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_reset; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_clock; // @[ClockGroup.scala 79:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_reset; // @[ClockGroup.scala 79:81]
  wire [29:0] dummyClockGroupSourceNode_io_covSum; // @[ClockGroup.scala 79:81]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_ready; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_valid; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_opcode; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_param; // @[SystemBus.scala 24:26]
  wire [3:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_size; // @[SystemBus.scala 24:26]
  wire [5:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_source; // @[SystemBus.scala 24:26]
  wire [31:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_address; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_bufferable; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_modifiable; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_readalloc; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_writealloc; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_privileged; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_secure; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_fetch; // @[SystemBus.scala 24:26]
  wire [7:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_mask; // @[SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_data; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_ready; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_valid; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_opcode; // @[SystemBus.scala 24:26]
  wire [3:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_size; // @[SystemBus.scala 24:26]
  wire [5:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_source; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_denied; // @[SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_data; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_corrupt; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size; // @[SystemBus.scala 24:26]
  wire [6:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source; // @[SystemBus.scala 24:26]
  wire [31:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_bufferable; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_modifiable; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_readalloc; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_writealloc; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_privileged; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_secure; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_fetch; // @[SystemBus.scala 24:26]
  wire [7:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask; // @[SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size; // @[SystemBus.scala 24:26]
  wire [6:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied; // @[SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param; // @[SystemBus.scala 24:26]
  wire [3:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size; // @[SystemBus.scala 24:26]
  wire [3:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source; // @[SystemBus.scala 24:26]
  wire [31:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_bufferable; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_modifiable; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_readalloc; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_writealloc; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_privileged; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_secure; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_fetch; // @[SystemBus.scala 24:26]
  wire [7:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask; // @[SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode; // @[SystemBus.scala 24:26]
  wire [3:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size; // @[SystemBus.scala 24:26]
  wire [3:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied; // @[SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param; // @[SystemBus.scala 24:26]
  wire [3:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size; // @[SystemBus.scala 24:26]
  wire [6:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source; // @[SystemBus.scala 24:26]
  wire [30:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address; // @[SystemBus.scala 24:26]
  wire [7:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask; // @[SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid; // @[SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode; // @[SystemBus.scala 24:26]
  wire [3:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size; // @[SystemBus.scala 24:26]
  wire [6:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied; // @[SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_fixedClockNode_out_1_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_fixedClockNode_out_1_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset; // @[SystemBus.scala 24:26]
  wire [29:0] subsystem_sbus_io_covSum; // @[SystemBus.scala 24:26]
  wire  subsystem_sbus_metaReset; // @[SystemBus.scala 24:26]
  wire  subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source; // @[PeripheryBus.scala 31:26]
  wire [30:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address; // @[PeripheryBus.scala 31:26]
  wire [7:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_fixedClockNode_out_clock; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_fixedClockNode_out_reset; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_bus_xing_in_a_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_bus_xing_in_a_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_pbus_auto_bus_xing_in_a_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_pbus_auto_bus_xing_in_a_bits_param; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_pbus_auto_bus_xing_in_a_bits_size; // @[PeripheryBus.scala 31:26]
  wire [6:0] subsystem_pbus_auto_bus_xing_in_a_bits_source; // @[PeripheryBus.scala 31:26]
  wire [30:0] subsystem_pbus_auto_bus_xing_in_a_bits_address; // @[PeripheryBus.scala 31:26]
  wire [7:0] subsystem_pbus_auto_bus_xing_in_a_bits_mask; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_pbus_auto_bus_xing_in_a_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_bus_xing_in_d_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_bus_xing_in_d_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_pbus_auto_bus_xing_in_d_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_pbus_auto_bus_xing_in_d_bits_size; // @[PeripheryBus.scala 31:26]
  wire [6:0] subsystem_pbus_auto_bus_xing_in_d_bits_source; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_bus_xing_in_d_bits_denied; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_pbus_auto_bus_xing_in_d_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_bus_xing_in_d_bits_corrupt; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_clock; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_reset; // @[PeripheryBus.scala 31:26]
  wire [29:0] subsystem_pbus_io_covSum; // @[PeripheryBus.scala 31:26]
  wire  subsystem_pbus_metaReset; // @[PeripheryBus.scala 31:26]
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_ready;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_valid;
  wire [7:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_id;
  wire [31:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_addr;
  wire [7:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_len;
  wire [2:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_size;
  wire [1:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_burst;
  wire [3:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_cache;
  wire [2:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_prot;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_ready;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_valid;
  wire [63:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_bits_data;
  wire [7:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_bits_strb;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_bits_last;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_ready;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_valid;
  wire [7:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_bits_id;
  wire [1:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_bits_resp;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_ready;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_valid;
  wire [7:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_id;
  wire [31:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_addr;
  wire [7:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_len;
  wire [2:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_size;
  wire [1:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_burst;
  wire [3:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_cache;
  wire [2:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_prot;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_ready;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_valid;
  wire [7:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_id;
  wire [63:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_data;
  wire [1:0] subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_resp;
  wire  subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_last;
  wire  subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock;
  wire  subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset;
  wire  subsystem_fbus_auto_bus_xing_out_a_ready;
  wire  subsystem_fbus_auto_bus_xing_out_a_valid;
  wire [2:0] subsystem_fbus_auto_bus_xing_out_a_bits_opcode;
  wire [2:0] subsystem_fbus_auto_bus_xing_out_a_bits_param;
  wire [3:0] subsystem_fbus_auto_bus_xing_out_a_bits_size;
  wire [3:0] subsystem_fbus_auto_bus_xing_out_a_bits_source;
  wire [31:0] subsystem_fbus_auto_bus_xing_out_a_bits_address;
  wire  subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_bufferable;
  wire  subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_modifiable;
  wire  subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_readalloc;
  wire  subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_writealloc;
  wire  subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_privileged;
  wire  subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_secure;
  wire  subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_fetch;
  wire [7:0] subsystem_fbus_auto_bus_xing_out_a_bits_mask;
  wire [63:0] subsystem_fbus_auto_bus_xing_out_a_bits_data;
  wire  subsystem_fbus_auto_bus_xing_out_d_ready;
  wire  subsystem_fbus_auto_bus_xing_out_d_valid;
  wire [2:0] subsystem_fbus_auto_bus_xing_out_d_bits_opcode;
  wire [3:0] subsystem_fbus_auto_bus_xing_out_d_bits_size;
  wire [3:0] subsystem_fbus_auto_bus_xing_out_d_bits_source;
  wire  subsystem_fbus_auto_bus_xing_out_d_bits_denied;
  wire [63:0] subsystem_fbus_auto_bus_xing_out_d_bits_data;
  wire  subsystem_fbus_auto_bus_xing_out_d_bits_corrupt;
  wire  subsystem_fbus_subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_clock;
  wire  subsystem_fbus_subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_reset;
  wire  subsystem_fbus_subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_clock;
  wire  subsystem_fbus_subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_reset;
  wire  subsystem_fbus_clockGroup_auto_in_member_subsystem_fbus_0_clock;
  wire  subsystem_fbus_clockGroup_auto_in_member_subsystem_fbus_0_reset;
  wire  subsystem_fbus_clockGroup_auto_out_clock;
  wire  subsystem_fbus_clockGroup_auto_out_reset;
  wire  subsystem_fbus_fixedClockNode_auto_in_clock;
  wire  subsystem_fbus_fixedClockNode_auto_in_reset;
  wire  subsystem_fbus_fixedClockNode_auto_out_clock;
  wire  subsystem_fbus_fixedClockNode_auto_out_reset;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_a_ready;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_a_valid;
  wire [2:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_opcode;
  wire [2:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_param;
  wire [3:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_size;
  wire [3:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_source;
  wire [31:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_address;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_bufferable;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_modifiable;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_readalloc;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_writealloc;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_privileged;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_secure;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_fetch;
  wire [7:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_mask;
  wire [63:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_data;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_d_ready;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_d_valid;
  wire [2:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_opcode;
  wire [3:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_size;
  wire [3:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_source;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_denied;
  wire [63:0] subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_data;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_corrupt;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_a_ready;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_a_valid;
  wire [2:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_opcode;
  wire [2:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_param;
  wire [3:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_size;
  wire [3:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_source;
  wire [31:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_address;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_bufferable;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_modifiable;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_readalloc;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_writealloc;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_privileged;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_secure;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_mask;
  wire [63:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_data;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_d_ready;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_d_valid;
  wire [2:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_opcode;
  wire [3:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_size;
  wire [3:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_source;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_denied;
  wire [63:0] subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_data;
  wire  subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_corrupt;
  wire  subsystem_fbus_buffer_clock; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_reset; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_a_ready; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] subsystem_fbus_buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] subsystem_fbus_buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] subsystem_fbus_buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28]
  wire [3:0] subsystem_fbus_buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28]
  wire [31:0] subsystem_fbus_buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_bufferable; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_modifiable; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_readalloc; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_writealloc; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_privileged; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_secure; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_fetch; // @[Buffer.scala 68:28]
  wire [7:0] subsystem_fbus_buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] subsystem_fbus_buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_d_ready; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] subsystem_fbus_buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] subsystem_fbus_buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28]
  wire [3:0] subsystem_fbus_buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] subsystem_fbus_buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_a_ready; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_a_valid; // @[Buffer.scala 68:28]
  wire [2:0] subsystem_fbus_buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28]
  wire [2:0] subsystem_fbus_buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28]
  wire [3:0] subsystem_fbus_buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28]
  wire [3:0] subsystem_fbus_buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28]
  wire [31:0] subsystem_fbus_buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_bufferable; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_modifiable; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_readalloc; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_writealloc; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_privileged; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_secure; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_fetch; // @[Buffer.scala 68:28]
  wire [7:0] subsystem_fbus_buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28]
  wire [63:0] subsystem_fbus_buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_d_ready; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_d_valid; // @[Buffer.scala 68:28]
  wire [2:0] subsystem_fbus_buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28]
  wire [3:0] subsystem_fbus_buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28]
  wire [3:0] subsystem_fbus_buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_d_bits_denied; // @[Buffer.scala 68:28]
  wire [63:0] subsystem_fbus_buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_buffer_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28]
  wire [29:0] subsystem_fbus_buffer_io_covSum; // @[Buffer.scala 68:28]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_clock; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_reset; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_ready; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_valid; // @[LazyModule.scala 432:27]
  wire [7:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_id; // @[LazyModule.scala 432:27]
  wire [31:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_addr; // @[LazyModule.scala 432:27]
  wire [7:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_len; // @[LazyModule.scala 432:27]
  wire [2:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_size; // @[LazyModule.scala 432:27]
  wire [1:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_burst; // @[LazyModule.scala 432:27]
  wire [3:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_cache; // @[LazyModule.scala 432:27]
  wire [2:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_prot; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_ready; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_valid; // @[LazyModule.scala 432:27]
  wire [63:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_bits_data; // @[LazyModule.scala 432:27]
  wire [7:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_bits_strb; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_bits_last; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_ready; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_valid; // @[LazyModule.scala 432:27]
  wire [7:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_bits_id; // @[LazyModule.scala 432:27]
  wire [1:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_bits_resp; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_ready; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_valid; // @[LazyModule.scala 432:27]
  wire [7:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_id; // @[LazyModule.scala 432:27]
  wire [31:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_addr; // @[LazyModule.scala 432:27]
  wire [7:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_len; // @[LazyModule.scala 432:27]
  wire [2:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_size; // @[LazyModule.scala 432:27]
  wire [1:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_burst; // @[LazyModule.scala 432:27]
  wire [3:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_cache; // @[LazyModule.scala 432:27]
  wire [2:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_prot; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_ready; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_valid; // @[LazyModule.scala 432:27]
  wire [7:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_id; // @[LazyModule.scala 432:27]
  wire [63:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_data; // @[LazyModule.scala 432:27]
  wire [1:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_resp; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_last; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_ready; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_valid; // @[LazyModule.scala 432:27]
  wire [2:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_opcode; // @[LazyModule.scala 432:27]
  wire [2:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_param; // @[LazyModule.scala 432:27]
  wire [3:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_size; // @[LazyModule.scala 432:27]
  wire [3:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_source; // @[LazyModule.scala 432:27]
  wire [31:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_address; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 432:27]
  wire [7:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_mask; // @[LazyModule.scala 432:27]
  wire [63:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_data; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_ready; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_valid; // @[LazyModule.scala 432:27]
  wire [2:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_opcode; // @[LazyModule.scala 432:27]
  wire [3:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_size; // @[LazyModule.scala 432:27]
  wire [3:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_source; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_denied; // @[LazyModule.scala 432:27]
  wire [63:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_data; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_corrupt; // @[LazyModule.scala 432:27]
  wire [29:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_io_covSum; // @[LazyModule.scala 432:27]
  wire  subsystem_fbus_coupler_from_port_named_slave_port_axi4_metaReset; // @[LazyModule.scala 432:27]
  wire  subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_source; // @[PeripheryBus.scala 31:26]
  wire [11:0] subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_address; // @[PeripheryBus.scala 31:26]
  wire [7:0] subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_mask; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_source; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_valid; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_bits_size; // @[PeripheryBus.scala 31:26]
  wire [11:0] subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_bits_source; // @[PeripheryBus.scala 31:26]
  wire [17:0] subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_bits_address; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_valid; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_bits_size; // @[PeripheryBus.scala 31:26]
  wire [11:0] subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_bits_source; // @[PeripheryBus.scala 31:26]
  wire [31:0] subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source; // @[PeripheryBus.scala 31:26]
  wire [16:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_valid; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_source; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_source; // @[PeripheryBus.scala 31:26]
  wire [25:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_address; // @[PeripheryBus.scala 31:26]
  wire [7:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_mask; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_source; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_source; // @[PeripheryBus.scala 31:26]
  wire [27:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_address; // @[PeripheryBus.scala 31:26]
  wire [7:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_mask; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_size; // @[PeripheryBus.scala 31:26]
  wire [10:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_source; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size; // @[PeripheryBus.scala 31:26]
  wire [6:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source; // @[PeripheryBus.scala 31:26]
  wire [30:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address; // @[PeripheryBus.scala 31:26]
  wire [7:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size; // @[PeripheryBus.scala 31:26]
  wire [6:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_fixedClockNode_out_0_clock; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_fixedClockNode_out_0_reset; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_a_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_a_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_bus_xing_in_a_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_bus_xing_in_a_bits_param; // @[PeripheryBus.scala 31:26]
  wire [3:0] subsystem_cbus_auto_bus_xing_in_a_bits_size; // @[PeripheryBus.scala 31:26]
  wire [6:0] subsystem_cbus_auto_bus_xing_in_a_bits_source; // @[PeripheryBus.scala 31:26]
  wire [30:0] subsystem_cbus_auto_bus_xing_in_a_bits_address; // @[PeripheryBus.scala 31:26]
  wire [7:0] subsystem_cbus_auto_bus_xing_in_a_bits_mask; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_bus_xing_in_a_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_d_ready; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_d_valid; // @[PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_bus_xing_in_d_bits_opcode; // @[PeripheryBus.scala 31:26]
  wire [3:0] subsystem_cbus_auto_bus_xing_in_d_bits_size; // @[PeripheryBus.scala 31:26]
  wire [6:0] subsystem_cbus_auto_bus_xing_in_d_bits_source; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_d_bits_denied; // @[PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_bus_xing_in_d_bits_data; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_d_bits_corrupt; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_clock; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_reset; // @[PeripheryBus.scala 31:26]
  wire [29:0] subsystem_cbus_io_covSum; // @[PeripheryBus.scala 31:26]
  wire  subsystem_cbus_metaReset; // @[PeripheryBus.scala 31:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid; // @[MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id; // @[MemoryBus.scala 25:26]
  wire [31:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr; // @[MemoryBus.scala 25:26]
  wire [7:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len; // @[MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size; // @[MemoryBus.scala 25:26]
  wire [1:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_lock; // @[MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_cache; // @[MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_prot; // @[MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_qos; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid; // @[MemoryBus.scala 25:26]
  wire [63:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data; // @[MemoryBus.scala 25:26]
  wire [7:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid; // @[MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id; // @[MemoryBus.scala 25:26]
  wire [1:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid; // @[MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id; // @[MemoryBus.scala 25:26]
  wire [31:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr; // @[MemoryBus.scala 25:26]
  wire [7:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len; // @[MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size; // @[MemoryBus.scala 25:26]
  wire [1:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_lock; // @[MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_cache; // @[MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_prot; // @[MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_qos; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid; // @[MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id; // @[MemoryBus.scala 25:26]
  wire [63:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data; // @[MemoryBus.scala 25:26]
  wire [1:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_ready; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_valid; // @[MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_bus_xing_in_a_bits_opcode; // @[MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_bus_xing_in_a_bits_size; // @[MemoryBus.scala 25:26]
  wire [8:0] subsystem_mbus_auto_bus_xing_in_a_bits_source; // @[MemoryBus.scala 25:26]
  wire [31:0] subsystem_mbus_auto_bus_xing_in_a_bits_address; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_bufferable; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_modifiable; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_readalloc; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_writealloc; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_privileged; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_secure; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_fetch; // @[MemoryBus.scala 25:26]
  wire [7:0] subsystem_mbus_auto_bus_xing_in_a_bits_mask; // @[MemoryBus.scala 25:26]
  wire [63:0] subsystem_mbus_auto_bus_xing_in_a_bits_data; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_d_ready; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_d_valid; // @[MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_bus_xing_in_d_bits_opcode; // @[MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_bus_xing_in_d_bits_size; // @[MemoryBus.scala 25:26]
  wire [8:0] subsystem_mbus_auto_bus_xing_in_d_bits_source; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_d_bits_denied; // @[MemoryBus.scala 25:26]
  wire [63:0] subsystem_mbus_auto_bus_xing_in_d_bits_data; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_d_bits_corrupt; // @[MemoryBus.scala 25:26]
  wire [29:0] subsystem_mbus_io_covSum; // @[MemoryBus.scala 25:26]
  wire  subsystem_mbus_metaReset; // @[MemoryBus.scala 25:26]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid; // @[BankedL2Params.scala 47:31]
  wire [2:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode; // @[BankedL2Params.scala 47:31]
  wire [2:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size; // @[BankedL2Params.scala 47:31]
  wire [8:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source; // @[BankedL2Params.scala 47:31]
  wire [31:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_bufferable; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_modifiable; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_readalloc; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_writealloc; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_privileged; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_secure; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_fetch; // @[BankedL2Params.scala 47:31]
  wire [7:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask; // @[BankedL2Params.scala 47:31]
  wire [63:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid; // @[BankedL2Params.scala 47:31]
  wire [2:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode; // @[BankedL2Params.scala 47:31]
  wire [2:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size; // @[BankedL2Params.scala 47:31]
  wire [8:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied; // @[BankedL2Params.scala 47:31]
  wire [63:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_ready; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_valid; // @[BankedL2Params.scala 47:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_opcode; // @[BankedL2Params.scala 47:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_size; // @[BankedL2Params.scala 47:31]
  wire [6:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_source; // @[BankedL2Params.scala 47:31]
  wire [31:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_address; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_bufferable; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_modifiable; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_readalloc; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_writealloc; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_privileged; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_secure; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_fetch; // @[BankedL2Params.scala 47:31]
  wire [7:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_mask; // @[BankedL2Params.scala 47:31]
  wire [63:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_data; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_d_ready; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_d_valid; // @[BankedL2Params.scala 47:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_opcode; // @[BankedL2Params.scala 47:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_size; // @[BankedL2Params.scala 47:31]
  wire [6:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_source; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_denied; // @[BankedL2Params.scala 47:31]
  wire [63:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_data; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_corrupt; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset; // @[BankedL2Params.scala 47:31]
  wire [29:0] subsystem_l2_wrapper_io_covSum; // @[BankedL2Params.scala 47:31]
  wire  subsystem_l2_wrapper_metaReset; // @[BankedL2Params.scala 47:31]
  wire  tile_prci_domain_auto_tile_reset_domain_cva6_tile_hartid_in; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_int_out_clock_xing_out_2_sync_0; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_int_out_clock_xing_out_1_sync_0; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_int_out_clock_xing_out_0_sync_0; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_int_in_clock_xing_in_2_sync_0; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_int_in_clock_xing_in_1_sync_0; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_int_in_clock_xing_in_0_sync_0; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_int_in_clock_xing_in_0_sync_1; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_ready; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_valid; // @[HasTiles.scala 252:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode; // @[HasTiles.scala 252:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param; // @[HasTiles.scala 252:38]
  wire [3:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size; // @[HasTiles.scala 252:38]
  wire [5:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source; // @[HasTiles.scala 252:38]
  wire [31:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_bufferable; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_modifiable; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_readalloc; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_writealloc; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_privileged; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_secure; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_fetch; // @[HasTiles.scala 252:38]
  wire [7:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask; // @[HasTiles.scala 252:38]
  wire [63:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_d_ready; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_d_valid; // @[HasTiles.scala 252:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_opcode; // @[HasTiles.scala 252:38]
  wire [3:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_size; // @[HasTiles.scala 252:38]
  wire [5:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_source; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_denied; // @[HasTiles.scala 252:38]
  wire [63:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_data; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_corrupt; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tap_clock_in_clock; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_auto_tap_clock_in_reset; // @[HasTiles.scala 252:38]
  wire [29:0] tile_prci_domain_io_covSum; // @[HasTiles.scala 252:38]
  wire  tile_prci_domain_metaReset; // @[HasTiles.scala 252:38]
  wire  plicDomainWrapper_auto_plic_int_in_0; // @[Plic.scala 359:39]
  wire  plicDomainWrapper_auto_plic_int_out_1_0; // @[Plic.scala 359:39]
  wire  plicDomainWrapper_auto_plic_int_out_0_0; // @[Plic.scala 359:39]
  wire  plicDomainWrapper_auto_plic_in_a_ready; // @[Plic.scala 359:39]
  wire  plicDomainWrapper_auto_plic_in_a_valid; // @[Plic.scala 359:39]
  wire [2:0] plicDomainWrapper_auto_plic_in_a_bits_opcode; // @[Plic.scala 359:39]
  wire [1:0] plicDomainWrapper_auto_plic_in_a_bits_size; // @[Plic.scala 359:39]
  wire [10:0] plicDomainWrapper_auto_plic_in_a_bits_source; // @[Plic.scala 359:39]
  wire [27:0] plicDomainWrapper_auto_plic_in_a_bits_address; // @[Plic.scala 359:39]
  wire [7:0] plicDomainWrapper_auto_plic_in_a_bits_mask; // @[Plic.scala 359:39]
  wire [63:0] plicDomainWrapper_auto_plic_in_a_bits_data; // @[Plic.scala 359:39]
  wire  plicDomainWrapper_auto_plic_in_d_ready; // @[Plic.scala 359:39]
  wire  plicDomainWrapper_auto_plic_in_d_valid; // @[Plic.scala 359:39]
  wire [2:0] plicDomainWrapper_auto_plic_in_d_bits_opcode; // @[Plic.scala 359:39]
  wire [1:0] plicDomainWrapper_auto_plic_in_d_bits_size; // @[Plic.scala 359:39]
  wire [10:0] plicDomainWrapper_auto_plic_in_d_bits_source; // @[Plic.scala 359:39]
  wire [63:0] plicDomainWrapper_auto_plic_in_d_bits_data; // @[Plic.scala 359:39]
  wire  plicDomainWrapper_auto_clock_in_clock; // @[Plic.scala 359:39]
  wire  plicDomainWrapper_auto_clock_in_reset; // @[Plic.scala 359:39]
  wire [29:0] plicDomainWrapper_io_covSum; // @[Plic.scala 359:39]
  wire  plicDomainWrapper_metaReset; // @[Plic.scala 359:39]
  wire  clint_clock; // @[CLINT.scala 109:27]
  wire  clint_reset; // @[CLINT.scala 109:27]
  wire  clint_auto_int_out_0; // @[CLINT.scala 109:27]
  wire  clint_auto_int_out_1; // @[CLINT.scala 109:27]
  wire  clint_auto_in_a_ready; // @[CLINT.scala 109:27]
  wire  clint_auto_in_a_valid; // @[CLINT.scala 109:27]
  wire [2:0] clint_auto_in_a_bits_opcode; // @[CLINT.scala 109:27]
  wire [1:0] clint_auto_in_a_bits_size; // @[CLINT.scala 109:27]
  wire [10:0] clint_auto_in_a_bits_source; // @[CLINT.scala 109:27]
  wire [25:0] clint_auto_in_a_bits_address; // @[CLINT.scala 109:27]
  wire [7:0] clint_auto_in_a_bits_mask; // @[CLINT.scala 109:27]
  wire [63:0] clint_auto_in_a_bits_data; // @[CLINT.scala 109:27]
  wire  clint_auto_in_d_ready; // @[CLINT.scala 109:27]
  wire  clint_auto_in_d_valid; // @[CLINT.scala 109:27]
  wire [2:0] clint_auto_in_d_bits_opcode; // @[CLINT.scala 109:27]
  wire [1:0] clint_auto_in_d_bits_size; // @[CLINT.scala 109:27]
  wire [10:0] clint_auto_in_d_bits_source; // @[CLINT.scala 109:27]
  wire [63:0] clint_auto_in_d_bits_data; // @[CLINT.scala 109:27]
  wire  clint_io_rtcTick; // @[CLINT.scala 109:27]
  wire [29:0] clint_io_covSum; // @[CLINT.scala 109:27]
  wire  xbar_auto_int_in_0; // @[Xbar.scala 30:26]
  wire  xbar_auto_int_out_0; // @[Xbar.scala 30:26]
  wire [29:0] xbar_io_covSum; // @[Xbar.scala 30:26]
  wire  xbar_1_auto_int_in_0; // @[Xbar.scala 30:26]
  wire  xbar_1_auto_int_out_0; // @[Xbar.scala 30:26]
  wire [29:0] xbar_1_io_covSum; // @[Xbar.scala 30:26]
  wire  xbar_2_auto_int_in_0; // @[Xbar.scala 30:26]
  wire  xbar_2_auto_int_out_0; // @[Xbar.scala 30:26]
  wire [29:0] xbar_2_io_covSum; // @[Xbar.scala 30:26]
  wire  tileHartIdNexusNode_auto_out; // @[HasTiles.scala 159:39]
  wire [29:0] tileHartIdNexusNode_io_covSum; // @[HasTiles.scala 159:39]
  wire  intsource_clock; // @[Crossing.scala 26:31]
  wire  intsource_reset; // @[Crossing.scala 26:31]
  wire  intsource_auto_in_0; // @[Crossing.scala 26:31]
  wire  intsource_auto_in_1; // @[Crossing.scala 26:31]
  wire  intsource_auto_out_sync_0; // @[Crossing.scala 26:31]
  wire  intsource_auto_out_sync_1; // @[Crossing.scala 26:31]
  wire [29:0] intsource_io_covSum; // @[Crossing.scala 26:31]
  wire  intsource_1_clock; // @[Crossing.scala 26:31]
  wire  intsource_1_reset; // @[Crossing.scala 26:31]
  wire  intsource_1_auto_in_0; // @[Crossing.scala 26:31]
  wire  intsource_1_auto_out_sync_0; // @[Crossing.scala 26:31]
  wire [29:0] intsource_1_io_covSum; // @[Crossing.scala 26:31]
  wire  intsource_2_clock; // @[Crossing.scala 26:31]
  wire  intsource_2_reset; // @[Crossing.scala 26:31]
  wire  intsource_2_auto_in_0; // @[Crossing.scala 26:31]
  wire  intsource_2_auto_out_sync_0; // @[Crossing.scala 26:31]
  wire [29:0] intsource_2_io_covSum; // @[Crossing.scala 26:31]
  wire  intsink_1_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_1_auto_out_0; // @[Crossing.scala 94:29]
  wire [29:0] intsink_1_io_covSum; // @[Crossing.scala 94:29]
  wire  intsink_2_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_2_auto_out_0; // @[Crossing.scala 94:29]
  wire [29:0] intsink_2_io_covSum; // @[Crossing.scala 94:29]
  wire  intsink_3_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_3_auto_out_0; // @[Crossing.scala 94:29]
  wire [29:0] intsink_3_io_covSum; // @[Crossing.scala 94:29]
  wire  bootROMDomainWrapper_auto_bootrom_in_a_ready; // @[BootROM.scala 70:42]
  wire  bootROMDomainWrapper_auto_bootrom_in_a_valid; // @[BootROM.scala 70:42]
  wire [1:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_size; // @[BootROM.scala 70:42]
  wire [10:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_source; // @[BootROM.scala 70:42]
  wire [16:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_address; // @[BootROM.scala 70:42]
  wire  bootROMDomainWrapper_auto_bootrom_in_d_ready; // @[BootROM.scala 70:42]
  wire  bootROMDomainWrapper_auto_bootrom_in_d_valid; // @[BootROM.scala 70:42]
  wire [1:0] bootROMDomainWrapper_auto_bootrom_in_d_bits_size; // @[BootROM.scala 70:42]
  wire [10:0] bootROMDomainWrapper_auto_bootrom_in_d_bits_source; // @[BootROM.scala 70:42]
  wire [63:0] bootROMDomainWrapper_auto_bootrom_in_d_bits_data; // @[BootROM.scala 70:42]
  wire [29:0] bootROMDomainWrapper_io_covSum; // @[BootROM.scala 70:42]
  wire  maskROM_clock; // @[MaskROM.scala 66:29]
  wire  maskROM_reset; // @[MaskROM.scala 66:29]
  wire  maskROM_auto_in_a_ready; // @[MaskROM.scala 66:29]
  wire  maskROM_auto_in_a_valid; // @[MaskROM.scala 66:29]
  wire [1:0] maskROM_auto_in_a_bits_size; // @[MaskROM.scala 66:29]
  wire [11:0] maskROM_auto_in_a_bits_source; // @[MaskROM.scala 66:29]
  wire [17:0] maskROM_auto_in_a_bits_address; // @[MaskROM.scala 66:29]
  wire  maskROM_auto_in_d_ready; // @[MaskROM.scala 66:29]
  wire  maskROM_auto_in_d_valid; // @[MaskROM.scala 66:29]
  wire [1:0] maskROM_auto_in_d_bits_size; // @[MaskROM.scala 66:29]
  wire [11:0] maskROM_auto_in_d_bits_source; // @[MaskROM.scala 66:29]
  wire [31:0] maskROM_auto_in_d_bits_data; // @[MaskROM.scala 66:29]
  wire [29:0] maskROM_io_covSum; // @[MaskROM.scala 66:29]
  wire  maskROM_metaReset; // @[MaskROM.scala 66:29]
  wire  uartClockDomainWrapper_auto_uart_0_int_xing_out_sync_0; // @[UART.scala 242:44]
  wire  uartClockDomainWrapper_auto_uart_0_control_xing_in_a_ready; // @[UART.scala 242:44]
  wire  uartClockDomainWrapper_auto_uart_0_control_xing_in_a_valid; // @[UART.scala 242:44]
  wire [2:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_opcode; // @[UART.scala 242:44]
  wire [1:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_size; // @[UART.scala 242:44]
  wire [10:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_source; // @[UART.scala 242:44]
  wire [30:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_address; // @[UART.scala 242:44]
  wire [7:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_mask; // @[UART.scala 242:44]
  wire [63:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_data; // @[UART.scala 242:44]
  wire  uartClockDomainWrapper_auto_uart_0_control_xing_in_d_ready; // @[UART.scala 242:44]
  wire  uartClockDomainWrapper_auto_uart_0_control_xing_in_d_valid; // @[UART.scala 242:44]
  wire [2:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_opcode; // @[UART.scala 242:44]
  wire [1:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_size; // @[UART.scala 242:44]
  wire [10:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_source; // @[UART.scala 242:44]
  wire [63:0] uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_data; // @[UART.scala 242:44]
  wire  uartClockDomainWrapper_auto_uart_0_io_out_txd; // @[UART.scala 242:44]
  wire  uartClockDomainWrapper_auto_uart_0_io_out_rxd; // @[UART.scala 242:44]
  wire  uartClockDomainWrapper_auto_clock_in_clock; // @[UART.scala 242:44]
  wire  uartClockDomainWrapper_auto_clock_in_reset; // @[UART.scala 242:44]
  wire [29:0] uartClockDomainWrapper_io_covSum; // @[UART.scala 242:44]
  wire  uartClockDomainWrapper_metaReset; // @[UART.scala 242:44]
  wire  intsink_4_auto_in_sync_0; // @[Crossing.scala 94:29]
  wire  intsink_4_auto_out_0; // @[Crossing.scala 94:29]
  wire [29:0] intsink_4_io_covSum; // @[Crossing.scala 94:29]
  wire  magic_clock; // @[Magic.scala 90:27]
  wire  magic_reset; // @[Magic.scala 90:27]
  wire  magic_auto_in_a_ready; // @[Magic.scala 90:27]
  wire  magic_auto_in_a_valid; // @[Magic.scala 90:27]
  wire [2:0] magic_auto_in_a_bits_opcode; // @[Magic.scala 90:27]
  wire [1:0] magic_auto_in_a_bits_size; // @[Magic.scala 90:27]
  wire [10:0] magic_auto_in_a_bits_source; // @[Magic.scala 90:27]
  wire [11:0] magic_auto_in_a_bits_address; // @[Magic.scala 90:27]
  wire [7:0] magic_auto_in_a_bits_mask; // @[Magic.scala 90:27]
  wire  magic_auto_in_d_ready; // @[Magic.scala 90:27]
  wire  magic_auto_in_d_valid; // @[Magic.scala 90:27]
  wire [2:0] magic_auto_in_d_bits_opcode; // @[Magic.scala 90:27]
  wire [1:0] magic_auto_in_d_bits_size; // @[Magic.scala 90:27]
  wire [10:0] magic_auto_in_d_bits_source; // @[Magic.scala 90:27]
  wire [63:0] magic_auto_in_d_bits_data; // @[Magic.scala 90:27]
  wire [29:0] magic_io_covSum; // @[Magic.scala 90:27]
  reg [6:0] int_rtc_tick_value; // @[Counter.scala 62:40]
  wire  int_rtc_tick_wrap_wrap = int_rtc_tick_value == 7'h63; // @[Counter.scala 74:24]
  wire [6:0] _int_rtc_tick_wrap_value_T_1 = int_rtc_tick_value + 7'h1; // @[Counter.scala 78:24]
  wire [29:0] StarshipASICTop_covSum;
  wire [29:0] subsystem_fbus_coupler_from_port_named_slave_port_axi4_sum;
  wire [29:0] ibus_int_bus_sum;
  wire [29:0] intsink_2_sum;
  wire [29:0] subsystem_fbus_buffer_sum;
  wire [29:0] subsystem_l2_wrapper_sum;
  wire [29:0] tile_prci_domain_sum;
  wire [29:0] maskROM_sum;
  wire [29:0] subsystem_sbus_sum;
  wire [29:0] subsystem_cbus_sum;
  wire [29:0] bootROMDomainWrapper_sum;
  wire [29:0] xbar_1_sum;
  wire [29:0] intsink_1_sum;
  wire [29:0] uartClockDomainWrapper_sum;
  wire [29:0] intsource_1_sum;
  wire [29:0] tileHartIdNexusNode_sum;
  wire [29:0] dummyClockGroupSourceNode_sum;
  wire [29:0] magic_sum;
  wire [29:0] subsystem_pbus_sum;
  wire [29:0] xbar_sum;
  wire [29:0] xbar_2_sum;
  wire [29:0] subsystem_mbus_sum;
  wire [29:0] plicDomainWrapper_sum;
  wire [29:0] intsource_sum;
  wire [29:0] intsink_4_sum;
  wire [29:0] clint_sum;
  wire [29:0] intsource_2_sum;
  wire [29:0] intsink_3_sum;
  IntXbar ibus_int_bus ( // @[InterruptBus.scala 14:27]
    .auto_int_in_0(ibus_int_bus_auto_int_in_0),
    .auto_int_out_0(ibus_int_bus_auto_int_out_0),
    .io_covSum(ibus_int_bus_io_covSum)
  );
  SimpleClockGroupSource dummyClockGroupSourceNode ( // @[ClockGroup.scala 79:81]
    .clock(dummyClockGroupSourceNode_clock),
    .reset(dummyClockGroupSourceNode_reset),
    .auto_out_member_subsystem_sbus_5_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_clock),
    .auto_out_member_subsystem_sbus_5_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_reset),
    .auto_out_member_subsystem_sbus_4_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_clock),
    .auto_out_member_subsystem_sbus_4_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_reset),
    .auto_out_member_subsystem_sbus_3_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_clock),
    .auto_out_member_subsystem_sbus_3_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_reset),
    .auto_out_member_subsystem_sbus_2_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_clock),
    .auto_out_member_subsystem_sbus_2_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_reset),
    .auto_out_member_subsystem_sbus_1_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_clock),
    .auto_out_member_subsystem_sbus_1_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_reset),
    .auto_out_member_subsystem_sbus_0_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_clock),
    .auto_out_member_subsystem_sbus_0_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_reset),
    .io_covSum(dummyClockGroupSourceNode_io_covSum)
  );
  SystemBus subsystem_sbus ( // @[SystemBus.scala 24:26]
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_ready(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_ready),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_valid(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_valid),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_opcode(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_opcode),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_param(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_param),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_size(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_size),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_source(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_source),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_address(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_address),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_bufferable(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_bufferable),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_modifiable(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_modifiable),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_readalloc(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_readalloc),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_writealloc(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_writealloc),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_privileged(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_privileged),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_secure(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_secure),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_fetch(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_fetch),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_mask(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_mask),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_data(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_data),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_ready(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_ready),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_valid(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_valid),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_opcode(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_opcode),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_size(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_size),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_source(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_source),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_denied(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_denied),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_data(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_data),
    .auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_corrupt(
      subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_corrupt),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_bufferable(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_bufferable),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_modifiable(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_modifiable),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_readalloc(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_readalloc),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_writealloc(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_writealloc),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_privileged(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_privileged),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_secure(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_secure),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_fetch(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_fetch),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_bufferable(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_bufferable),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_modifiable(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_modifiable),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_readalloc(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_readalloc),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_writealloc(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_writealloc),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_privileged(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_privileged),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_secure(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_secure),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_fetch(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_fetch),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data),
    .auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt(
      subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt),
    .auto_fixedClockNode_out_1_clock(subsystem_sbus_auto_fixedClockNode_out_1_clock),
    .auto_fixedClockNode_out_1_reset(subsystem_sbus_auto_fixedClockNode_out_1_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset),
    .auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock),
    .auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset),
    .auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock),
    .auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset),
    .auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock),
    .auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset),
    .auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock),
    .auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset),
    .auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock),
    .auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset),
    .io_covSum(subsystem_sbus_io_covSum),
    .metaReset(subsystem_sbus_metaReset)
  );
  PeripheryBus subsystem_pbus ( // @[PeripheryBus.scala 31:26]
    .auto_coupler_to_device_named_uart_0_control_xing_out_a_ready(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_ready),
    .auto_coupler_to_device_named_uart_0_control_xing_out_a_valid(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_valid),
    .auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode),
    .auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size),
    .auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source),
    .auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address),
    .auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask),
    .auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data),
    .auto_coupler_to_device_named_uart_0_control_xing_out_d_ready(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_ready),
    .auto_coupler_to_device_named_uart_0_control_xing_out_d_valid(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_valid),
    .auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode),
    .auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size),
    .auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source),
    .auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data(
      subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data),
    .auto_fixedClockNode_out_clock(subsystem_pbus_auto_fixedClockNode_out_clock),
    .auto_fixedClockNode_out_reset(subsystem_pbus_auto_fixedClockNode_out_reset),
    .auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock(
      subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock),
    .auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset(
      subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset),
    .auto_bus_xing_in_a_ready(subsystem_pbus_auto_bus_xing_in_a_ready),
    .auto_bus_xing_in_a_valid(subsystem_pbus_auto_bus_xing_in_a_valid),
    .auto_bus_xing_in_a_bits_opcode(subsystem_pbus_auto_bus_xing_in_a_bits_opcode),
    .auto_bus_xing_in_a_bits_param(subsystem_pbus_auto_bus_xing_in_a_bits_param),
    .auto_bus_xing_in_a_bits_size(subsystem_pbus_auto_bus_xing_in_a_bits_size),
    .auto_bus_xing_in_a_bits_source(subsystem_pbus_auto_bus_xing_in_a_bits_source),
    .auto_bus_xing_in_a_bits_address(subsystem_pbus_auto_bus_xing_in_a_bits_address),
    .auto_bus_xing_in_a_bits_mask(subsystem_pbus_auto_bus_xing_in_a_bits_mask),
    .auto_bus_xing_in_a_bits_data(subsystem_pbus_auto_bus_xing_in_a_bits_data),
    .auto_bus_xing_in_d_ready(subsystem_pbus_auto_bus_xing_in_d_ready),
    .auto_bus_xing_in_d_valid(subsystem_pbus_auto_bus_xing_in_d_valid),
    .auto_bus_xing_in_d_bits_opcode(subsystem_pbus_auto_bus_xing_in_d_bits_opcode),
    .auto_bus_xing_in_d_bits_size(subsystem_pbus_auto_bus_xing_in_d_bits_size),
    .auto_bus_xing_in_d_bits_source(subsystem_pbus_auto_bus_xing_in_d_bits_source),
    .auto_bus_xing_in_d_bits_denied(subsystem_pbus_auto_bus_xing_in_d_bits_denied),
    .auto_bus_xing_in_d_bits_data(subsystem_pbus_auto_bus_xing_in_d_bits_data),
    .auto_bus_xing_in_d_bits_corrupt(subsystem_pbus_auto_bus_xing_in_d_bits_corrupt),
    .clock(subsystem_pbus_clock),
    .reset(subsystem_pbus_reset),
    .io_covSum(subsystem_pbus_io_covSum),
    .metaReset(subsystem_pbus_metaReset)
  );
  TLBuffer_2 subsystem_fbus_buffer ( // @[Buffer.scala 68:28]
    .clock(subsystem_fbus_buffer_clock),
    .reset(subsystem_fbus_buffer_reset),
    .auto_in_a_ready(subsystem_fbus_buffer_auto_in_a_ready),
    .auto_in_a_valid(subsystem_fbus_buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(subsystem_fbus_buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(subsystem_fbus_buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(subsystem_fbus_buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(subsystem_fbus_buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(subsystem_fbus_buffer_auto_in_a_bits_address),
    .auto_in_a_bits_user_amba_prot_bufferable(subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_bufferable),
    .auto_in_a_bits_user_amba_prot_modifiable(subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_modifiable),
    .auto_in_a_bits_user_amba_prot_readalloc(subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_readalloc),
    .auto_in_a_bits_user_amba_prot_writealloc(subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_writealloc),
    .auto_in_a_bits_user_amba_prot_privileged(subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_privileged),
    .auto_in_a_bits_user_amba_prot_secure(subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_secure),
    .auto_in_a_bits_user_amba_prot_fetch(subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_fetch),
    .auto_in_a_bits_mask(subsystem_fbus_buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(subsystem_fbus_buffer_auto_in_a_bits_data),
    .auto_in_d_ready(subsystem_fbus_buffer_auto_in_d_ready),
    .auto_in_d_valid(subsystem_fbus_buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(subsystem_fbus_buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(subsystem_fbus_buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(subsystem_fbus_buffer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(subsystem_fbus_buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(subsystem_fbus_buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(subsystem_fbus_buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(subsystem_fbus_buffer_auto_out_a_ready),
    .auto_out_a_valid(subsystem_fbus_buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(subsystem_fbus_buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(subsystem_fbus_buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(subsystem_fbus_buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(subsystem_fbus_buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(subsystem_fbus_buffer_auto_out_a_bits_address),
    .auto_out_a_bits_user_amba_prot_bufferable(subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_bufferable),
    .auto_out_a_bits_user_amba_prot_modifiable(subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_modifiable),
    .auto_out_a_bits_user_amba_prot_readalloc(subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_readalloc),
    .auto_out_a_bits_user_amba_prot_writealloc(subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_writealloc),
    .auto_out_a_bits_user_amba_prot_privileged(subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_privileged),
    .auto_out_a_bits_user_amba_prot_secure(subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_secure),
    .auto_out_a_bits_user_amba_prot_fetch(subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_fetch),
    .auto_out_a_bits_mask(subsystem_fbus_buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(subsystem_fbus_buffer_auto_out_a_bits_data),
    .auto_out_d_ready(subsystem_fbus_buffer_auto_out_d_ready),
    .auto_out_d_valid(subsystem_fbus_buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(subsystem_fbus_buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(subsystem_fbus_buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(subsystem_fbus_buffer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(subsystem_fbus_buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(subsystem_fbus_buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(subsystem_fbus_buffer_auto_out_d_bits_corrupt),
    .io_covSum(subsystem_fbus_buffer_io_covSum)
  );
  TLInterconnectCoupler_5 subsystem_fbus_coupler_from_port_named_slave_port_axi4 ( // @[LazyModule.scala 432:27]
    .clock(subsystem_fbus_coupler_from_port_named_slave_port_axi4_clock),
    .reset(subsystem_fbus_coupler_from_port_named_slave_port_axi4_reset),
    .auto_axi4index_in_aw_ready(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_ready),
    .auto_axi4index_in_aw_valid(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_valid),
    .auto_axi4index_in_aw_bits_id(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_id),
    .auto_axi4index_in_aw_bits_addr(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_addr),
    .auto_axi4index_in_aw_bits_len(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_len)
      ,
    .auto_axi4index_in_aw_bits_size(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_size),
    .auto_axi4index_in_aw_bits_burst(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_burst),
    .auto_axi4index_in_aw_bits_cache(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_cache),
    .auto_axi4index_in_aw_bits_prot(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_prot),
    .auto_axi4index_in_w_ready(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_ready),
    .auto_axi4index_in_w_valid(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_valid),
    .auto_axi4index_in_w_bits_data(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_bits_data)
      ,
    .auto_axi4index_in_w_bits_strb(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_bits_strb)
      ,
    .auto_axi4index_in_w_bits_last(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_bits_last)
      ,
    .auto_axi4index_in_b_ready(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_ready),
    .auto_axi4index_in_b_valid(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_valid),
    .auto_axi4index_in_b_bits_id(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_bits_id),
    .auto_axi4index_in_b_bits_resp(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_bits_resp)
      ,
    .auto_axi4index_in_ar_ready(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_ready),
    .auto_axi4index_in_ar_valid(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_valid),
    .auto_axi4index_in_ar_bits_id(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_id),
    .auto_axi4index_in_ar_bits_addr(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_addr),
    .auto_axi4index_in_ar_bits_len(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_len)
      ,
    .auto_axi4index_in_ar_bits_size(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_size),
    .auto_axi4index_in_ar_bits_burst(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_burst),
    .auto_axi4index_in_ar_bits_cache(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_cache),
    .auto_axi4index_in_ar_bits_prot(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_prot),
    .auto_axi4index_in_r_ready(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_ready),
    .auto_axi4index_in_r_valid(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_valid),
    .auto_axi4index_in_r_bits_id(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_id),
    .auto_axi4index_in_r_bits_data(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_data)
      ,
    .auto_axi4index_in_r_bits_resp(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_resp)
      ,
    .auto_axi4index_in_r_bits_last(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_last)
      ,
    .auto_tl_out_a_ready(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_ready),
    .auto_tl_out_a_valid(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_valid),
    .auto_tl_out_a_bits_opcode(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_opcode),
    .auto_tl_out_a_bits_param(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_param),
    .auto_tl_out_a_bits_size(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_size),
    .auto_tl_out_a_bits_source(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_source),
    .auto_tl_out_a_bits_address(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_address),
    .auto_tl_out_a_bits_user_amba_prot_bufferable(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_bufferable),
    .auto_tl_out_a_bits_user_amba_prot_modifiable(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_modifiable),
    .auto_tl_out_a_bits_user_amba_prot_readalloc(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_readalloc),
    .auto_tl_out_a_bits_user_amba_prot_writealloc(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_writealloc),
    .auto_tl_out_a_bits_user_amba_prot_privileged(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_privileged),
    .auto_tl_out_a_bits_user_amba_prot_secure(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_secure),
    .auto_tl_out_a_bits_user_amba_prot_fetch(
      subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_fetch),
    .auto_tl_out_a_bits_mask(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_mask),
    .auto_tl_out_a_bits_data(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_data),
    .auto_tl_out_d_ready(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_ready),
    .auto_tl_out_d_valid(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_valid),
    .auto_tl_out_d_bits_opcode(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_opcode),
    .auto_tl_out_d_bits_size(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_size),
    .auto_tl_out_d_bits_source(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_source),
    .auto_tl_out_d_bits_denied(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_denied),
    .auto_tl_out_d_bits_data(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_data),
    .auto_tl_out_d_bits_corrupt(subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_corrupt),
    .io_covSum(subsystem_fbus_coupler_from_port_named_slave_port_axi4_io_covSum),
    .metaReset(subsystem_fbus_coupler_from_port_named_slave_port_axi4_metaReset)
  );
  PeripheryBus_1 subsystem_cbus ( // @[PeripheryBus.scala 31:26]
    .auto_coupler_to_magic_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_ready),
    .auto_coupler_to_magic_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_valid),
    .auto_coupler_to_magic_fragmenter_out_a_bits_opcode(
      subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_opcode),
    .auto_coupler_to_magic_fragmenter_out_a_bits_size(subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_size),
    .auto_coupler_to_magic_fragmenter_out_a_bits_source(
      subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_source),
    .auto_coupler_to_magic_fragmenter_out_a_bits_address(
      subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_address),
    .auto_coupler_to_magic_fragmenter_out_a_bits_mask(subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_mask),
    .auto_coupler_to_magic_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_ready),
    .auto_coupler_to_magic_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_valid),
    .auto_coupler_to_magic_fragmenter_out_d_bits_opcode(
      subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_opcode),
    .auto_coupler_to_magic_fragmenter_out_d_bits_size(subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_size),
    .auto_coupler_to_magic_fragmenter_out_d_bits_source(
      subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_source),
    .auto_coupler_to_magic_fragmenter_out_d_bits_data(subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_data),
    .auto_coupler_to_MaskROM_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_ready),
    .auto_coupler_to_MaskROM_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_valid),
    .auto_coupler_to_MaskROM_fragmenter_out_a_bits_size(
      subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_bits_size),
    .auto_coupler_to_MaskROM_fragmenter_out_a_bits_source(
      subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_bits_source),
    .auto_coupler_to_MaskROM_fragmenter_out_a_bits_address(
      subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_bits_address),
    .auto_coupler_to_MaskROM_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_ready),
    .auto_coupler_to_MaskROM_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_valid),
    .auto_coupler_to_MaskROM_fragmenter_out_d_bits_size(
      subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_bits_size),
    .auto_coupler_to_MaskROM_fragmenter_out_d_bits_source(
      subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_bits_source),
    .auto_coupler_to_MaskROM_fragmenter_out_d_bits_data(
      subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_bits_data),
    .auto_coupler_to_bootrom_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_ready),
    .auto_coupler_to_bootrom_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid),
    .auto_coupler_to_bootrom_fragmenter_out_a_bits_size(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size),
    .auto_coupler_to_bootrom_fragmenter_out_a_bits_source(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source),
    .auto_coupler_to_bootrom_fragmenter_out_a_bits_address(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address),
    .auto_coupler_to_bootrom_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready),
    .auto_coupler_to_bootrom_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_valid),
    .auto_coupler_to_bootrom_fragmenter_out_d_bits_size(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_size),
    .auto_coupler_to_bootrom_fragmenter_out_d_bits_source(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_source),
    .auto_coupler_to_bootrom_fragmenter_out_d_bits_data(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_data),
    .auto_coupler_to_clint_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_ready),
    .auto_coupler_to_clint_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_valid),
    .auto_coupler_to_clint_fragmenter_out_a_bits_opcode(
      subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_opcode),
    .auto_coupler_to_clint_fragmenter_out_a_bits_size(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_size),
    .auto_coupler_to_clint_fragmenter_out_a_bits_source(
      subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_source),
    .auto_coupler_to_clint_fragmenter_out_a_bits_address(
      subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_address),
    .auto_coupler_to_clint_fragmenter_out_a_bits_mask(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_mask),
    .auto_coupler_to_clint_fragmenter_out_a_bits_data(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_data),
    .auto_coupler_to_clint_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_ready),
    .auto_coupler_to_clint_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_valid),
    .auto_coupler_to_clint_fragmenter_out_d_bits_opcode(
      subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_opcode),
    .auto_coupler_to_clint_fragmenter_out_d_bits_size(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_size),
    .auto_coupler_to_clint_fragmenter_out_d_bits_source(
      subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_source),
    .auto_coupler_to_clint_fragmenter_out_d_bits_data(subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_data),
    .auto_coupler_to_plic_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_ready),
    .auto_coupler_to_plic_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_valid),
    .auto_coupler_to_plic_fragmenter_out_a_bits_opcode(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_opcode)
      ,
    .auto_coupler_to_plic_fragmenter_out_a_bits_size(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_size),
    .auto_coupler_to_plic_fragmenter_out_a_bits_source(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_source)
      ,
    .auto_coupler_to_plic_fragmenter_out_a_bits_address(
      subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_address),
    .auto_coupler_to_plic_fragmenter_out_a_bits_mask(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_mask),
    .auto_coupler_to_plic_fragmenter_out_a_bits_data(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_data),
    .auto_coupler_to_plic_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_ready),
    .auto_coupler_to_plic_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_valid),
    .auto_coupler_to_plic_fragmenter_out_d_bits_opcode(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_opcode)
      ,
    .auto_coupler_to_plic_fragmenter_out_d_bits_size(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_size),
    .auto_coupler_to_plic_fragmenter_out_d_bits_source(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_source)
      ,
    .auto_coupler_to_plic_fragmenter_out_d_bits_data(subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_data),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data),
    .auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt(
      subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt),
    .auto_fixedClockNode_out_0_clock(subsystem_cbus_auto_fixedClockNode_out_0_clock),
    .auto_fixedClockNode_out_0_reset(subsystem_cbus_auto_fixedClockNode_out_0_reset),
    .auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock),
    .auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset),
    .auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock),
    .auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset),
    .auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock),
    .auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset),
    .auto_bus_xing_in_a_ready(subsystem_cbus_auto_bus_xing_in_a_ready),
    .auto_bus_xing_in_a_valid(subsystem_cbus_auto_bus_xing_in_a_valid),
    .auto_bus_xing_in_a_bits_opcode(subsystem_cbus_auto_bus_xing_in_a_bits_opcode),
    .auto_bus_xing_in_a_bits_param(subsystem_cbus_auto_bus_xing_in_a_bits_param),
    .auto_bus_xing_in_a_bits_size(subsystem_cbus_auto_bus_xing_in_a_bits_size),
    .auto_bus_xing_in_a_bits_source(subsystem_cbus_auto_bus_xing_in_a_bits_source),
    .auto_bus_xing_in_a_bits_address(subsystem_cbus_auto_bus_xing_in_a_bits_address),
    .auto_bus_xing_in_a_bits_mask(subsystem_cbus_auto_bus_xing_in_a_bits_mask),
    .auto_bus_xing_in_a_bits_data(subsystem_cbus_auto_bus_xing_in_a_bits_data),
    .auto_bus_xing_in_d_ready(subsystem_cbus_auto_bus_xing_in_d_ready),
    .auto_bus_xing_in_d_valid(subsystem_cbus_auto_bus_xing_in_d_valid),
    .auto_bus_xing_in_d_bits_opcode(subsystem_cbus_auto_bus_xing_in_d_bits_opcode),
    .auto_bus_xing_in_d_bits_size(subsystem_cbus_auto_bus_xing_in_d_bits_size),
    .auto_bus_xing_in_d_bits_source(subsystem_cbus_auto_bus_xing_in_d_bits_source),
    .auto_bus_xing_in_d_bits_denied(subsystem_cbus_auto_bus_xing_in_d_bits_denied),
    .auto_bus_xing_in_d_bits_data(subsystem_cbus_auto_bus_xing_in_d_bits_data),
    .auto_bus_xing_in_d_bits_corrupt(subsystem_cbus_auto_bus_xing_in_d_bits_corrupt),
    .clock(subsystem_cbus_clock),
    .reset(subsystem_cbus_reset),
    .io_covSum(subsystem_cbus_io_covSum),
    .metaReset(subsystem_cbus_metaReset)
  );
  MemoryBus subsystem_mbus ( // @[MemoryBus.scala 25:26]
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_lock(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_lock),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_cache(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_cache),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_prot(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_prot),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_qos(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_qos),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_lock(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_lock),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_cache(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_cache),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_prot(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_prot),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_qos(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_qos),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last),
    .auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock(
      subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock),
    .auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset(
      subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset),
    .auto_bus_xing_in_a_ready(subsystem_mbus_auto_bus_xing_in_a_ready),
    .auto_bus_xing_in_a_valid(subsystem_mbus_auto_bus_xing_in_a_valid),
    .auto_bus_xing_in_a_bits_opcode(subsystem_mbus_auto_bus_xing_in_a_bits_opcode),
    .auto_bus_xing_in_a_bits_size(subsystem_mbus_auto_bus_xing_in_a_bits_size),
    .auto_bus_xing_in_a_bits_source(subsystem_mbus_auto_bus_xing_in_a_bits_source),
    .auto_bus_xing_in_a_bits_address(subsystem_mbus_auto_bus_xing_in_a_bits_address),
    .auto_bus_xing_in_a_bits_user_amba_prot_bufferable(subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_bufferable)
      ,
    .auto_bus_xing_in_a_bits_user_amba_prot_modifiable(subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_modifiable)
      ,
    .auto_bus_xing_in_a_bits_user_amba_prot_readalloc(subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_readalloc),
    .auto_bus_xing_in_a_bits_user_amba_prot_writealloc(subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_writealloc)
      ,
    .auto_bus_xing_in_a_bits_user_amba_prot_privileged(subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_privileged)
      ,
    .auto_bus_xing_in_a_bits_user_amba_prot_secure(subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_secure),
    .auto_bus_xing_in_a_bits_user_amba_prot_fetch(subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_fetch),
    .auto_bus_xing_in_a_bits_mask(subsystem_mbus_auto_bus_xing_in_a_bits_mask),
    .auto_bus_xing_in_a_bits_data(subsystem_mbus_auto_bus_xing_in_a_bits_data),
    .auto_bus_xing_in_d_ready(subsystem_mbus_auto_bus_xing_in_d_ready),
    .auto_bus_xing_in_d_valid(subsystem_mbus_auto_bus_xing_in_d_valid),
    .auto_bus_xing_in_d_bits_opcode(subsystem_mbus_auto_bus_xing_in_d_bits_opcode),
    .auto_bus_xing_in_d_bits_size(subsystem_mbus_auto_bus_xing_in_d_bits_size),
    .auto_bus_xing_in_d_bits_source(subsystem_mbus_auto_bus_xing_in_d_bits_source),
    .auto_bus_xing_in_d_bits_denied(subsystem_mbus_auto_bus_xing_in_d_bits_denied),
    .auto_bus_xing_in_d_bits_data(subsystem_mbus_auto_bus_xing_in_d_bits_data),
    .auto_bus_xing_in_d_bits_corrupt(subsystem_mbus_auto_bus_xing_in_d_bits_corrupt),
    .io_covSum(subsystem_mbus_io_covSum),
    .metaReset(subsystem_mbus_metaReset)
  );
  CoherenceManagerWrapper subsystem_l2_wrapper ( // @[BankedL2Params.scala 47:31]
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_bufferable(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_bufferable),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_modifiable(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_modifiable),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_readalloc(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_readalloc),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_writealloc(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_writealloc),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_privileged(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_privileged),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_secure(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_secure),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_fetch(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_fetch),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt),
    .auto_coherent_jbar_in_a_ready(subsystem_l2_wrapper_auto_coherent_jbar_in_a_ready),
    .auto_coherent_jbar_in_a_valid(subsystem_l2_wrapper_auto_coherent_jbar_in_a_valid),
    .auto_coherent_jbar_in_a_bits_opcode(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_opcode),
    .auto_coherent_jbar_in_a_bits_size(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_size),
    .auto_coherent_jbar_in_a_bits_source(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_source),
    .auto_coherent_jbar_in_a_bits_address(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_address),
    .auto_coherent_jbar_in_a_bits_user_amba_prot_bufferable(
      subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_bufferable),
    .auto_coherent_jbar_in_a_bits_user_amba_prot_modifiable(
      subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_modifiable),
    .auto_coherent_jbar_in_a_bits_user_amba_prot_readalloc(
      subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_readalloc),
    .auto_coherent_jbar_in_a_bits_user_amba_prot_writealloc(
      subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_writealloc),
    .auto_coherent_jbar_in_a_bits_user_amba_prot_privileged(
      subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_privileged),
    .auto_coherent_jbar_in_a_bits_user_amba_prot_secure(
      subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_secure),
    .auto_coherent_jbar_in_a_bits_user_amba_prot_fetch(
      subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_fetch),
    .auto_coherent_jbar_in_a_bits_mask(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_mask),
    .auto_coherent_jbar_in_a_bits_data(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_data),
    .auto_coherent_jbar_in_d_ready(subsystem_l2_wrapper_auto_coherent_jbar_in_d_ready),
    .auto_coherent_jbar_in_d_valid(subsystem_l2_wrapper_auto_coherent_jbar_in_d_valid),
    .auto_coherent_jbar_in_d_bits_opcode(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_opcode),
    .auto_coherent_jbar_in_d_bits_size(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_size),
    .auto_coherent_jbar_in_d_bits_source(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_source),
    .auto_coherent_jbar_in_d_bits_denied(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_denied),
    .auto_coherent_jbar_in_d_bits_data(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_data),
    .auto_coherent_jbar_in_d_bits_corrupt(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_corrupt),
    .auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock),
    .auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset),
    .auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock),
    .auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset),
    .auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock),
    .auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset),
    .io_covSum(subsystem_l2_wrapper_io_covSum),
    .metaReset(subsystem_l2_wrapper_metaReset)
  );
  TilePRCIDomain tile_prci_domain ( // @[HasTiles.scala 252:38]
    .auto_tile_reset_domain_cva6_tile_hartid_in(tile_prci_domain_auto_tile_reset_domain_cva6_tile_hartid_in),
    .auto_int_out_clock_xing_out_2_sync_0(tile_prci_domain_auto_int_out_clock_xing_out_2_sync_0),
    .auto_int_out_clock_xing_out_1_sync_0(tile_prci_domain_auto_int_out_clock_xing_out_1_sync_0),
    .auto_int_out_clock_xing_out_0_sync_0(tile_prci_domain_auto_int_out_clock_xing_out_0_sync_0),
    .auto_int_in_clock_xing_in_2_sync_0(tile_prci_domain_auto_int_in_clock_xing_in_2_sync_0),
    .auto_int_in_clock_xing_in_1_sync_0(tile_prci_domain_auto_int_in_clock_xing_in_1_sync_0),
    .auto_int_in_clock_xing_in_0_sync_0(tile_prci_domain_auto_int_in_clock_xing_in_0_sync_0),
    .auto_int_in_clock_xing_in_0_sync_1(tile_prci_domain_auto_int_in_clock_xing_in_0_sync_1),
    .auto_tl_master_clock_xing_out_a_ready(tile_prci_domain_auto_tl_master_clock_xing_out_a_ready),
    .auto_tl_master_clock_xing_out_a_valid(tile_prci_domain_auto_tl_master_clock_xing_out_a_valid),
    .auto_tl_master_clock_xing_out_a_bits_opcode(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode),
    .auto_tl_master_clock_xing_out_a_bits_param(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param),
    .auto_tl_master_clock_xing_out_a_bits_size(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size),
    .auto_tl_master_clock_xing_out_a_bits_source(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source),
    .auto_tl_master_clock_xing_out_a_bits_address(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address),
    .auto_tl_master_clock_xing_out_a_bits_user_amba_prot_bufferable(
      tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_bufferable),
    .auto_tl_master_clock_xing_out_a_bits_user_amba_prot_modifiable(
      tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_modifiable),
    .auto_tl_master_clock_xing_out_a_bits_user_amba_prot_readalloc(
      tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_readalloc),
    .auto_tl_master_clock_xing_out_a_bits_user_amba_prot_writealloc(
      tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_writealloc),
    .auto_tl_master_clock_xing_out_a_bits_user_amba_prot_privileged(
      tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_privileged),
    .auto_tl_master_clock_xing_out_a_bits_user_amba_prot_secure(
      tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_secure),
    .auto_tl_master_clock_xing_out_a_bits_user_amba_prot_fetch(
      tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_fetch),
    .auto_tl_master_clock_xing_out_a_bits_mask(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask),
    .auto_tl_master_clock_xing_out_a_bits_data(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data),
    .auto_tl_master_clock_xing_out_d_ready(tile_prci_domain_auto_tl_master_clock_xing_out_d_ready),
    .auto_tl_master_clock_xing_out_d_valid(tile_prci_domain_auto_tl_master_clock_xing_out_d_valid),
    .auto_tl_master_clock_xing_out_d_bits_opcode(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_opcode),
    .auto_tl_master_clock_xing_out_d_bits_size(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_size),
    .auto_tl_master_clock_xing_out_d_bits_source(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_source),
    .auto_tl_master_clock_xing_out_d_bits_denied(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_denied),
    .auto_tl_master_clock_xing_out_d_bits_data(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_data),
    .auto_tl_master_clock_xing_out_d_bits_corrupt(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_corrupt),
    .auto_tap_clock_in_clock(tile_prci_domain_auto_tap_clock_in_clock),
    .auto_tap_clock_in_reset(tile_prci_domain_auto_tap_clock_in_reset),
    .io_covSum(tile_prci_domain_io_covSum),
    .metaReset(tile_prci_domain_metaReset)
  );
  ClockSinkDomain plicDomainWrapper ( // @[Plic.scala 359:39]
    .auto_plic_int_in_0(plicDomainWrapper_auto_plic_int_in_0),
    .auto_plic_int_out_1_0(plicDomainWrapper_auto_plic_int_out_1_0),
    .auto_plic_int_out_0_0(plicDomainWrapper_auto_plic_int_out_0_0),
    .auto_plic_in_a_ready(plicDomainWrapper_auto_plic_in_a_ready),
    .auto_plic_in_a_valid(plicDomainWrapper_auto_plic_in_a_valid),
    .auto_plic_in_a_bits_opcode(plicDomainWrapper_auto_plic_in_a_bits_opcode),
    .auto_plic_in_a_bits_size(plicDomainWrapper_auto_plic_in_a_bits_size),
    .auto_plic_in_a_bits_source(plicDomainWrapper_auto_plic_in_a_bits_source),
    .auto_plic_in_a_bits_address(plicDomainWrapper_auto_plic_in_a_bits_address),
    .auto_plic_in_a_bits_mask(plicDomainWrapper_auto_plic_in_a_bits_mask),
    .auto_plic_in_a_bits_data(plicDomainWrapper_auto_plic_in_a_bits_data),
    .auto_plic_in_d_ready(plicDomainWrapper_auto_plic_in_d_ready),
    .auto_plic_in_d_valid(plicDomainWrapper_auto_plic_in_d_valid),
    .auto_plic_in_d_bits_opcode(plicDomainWrapper_auto_plic_in_d_bits_opcode),
    .auto_plic_in_d_bits_size(plicDomainWrapper_auto_plic_in_d_bits_size),
    .auto_plic_in_d_bits_source(plicDomainWrapper_auto_plic_in_d_bits_source),
    .auto_plic_in_d_bits_data(plicDomainWrapper_auto_plic_in_d_bits_data),
    .auto_clock_in_clock(plicDomainWrapper_auto_clock_in_clock),
    .auto_clock_in_reset(plicDomainWrapper_auto_clock_in_reset),
    .io_covSum(plicDomainWrapper_io_covSum),
    .metaReset(plicDomainWrapper_metaReset)
  );
  CLINT clint ( // @[CLINT.scala 109:27]
    .clock(clint_clock),
    .reset(clint_reset),
    .auto_int_out_0(clint_auto_int_out_0),
    .auto_int_out_1(clint_auto_int_out_1),
    .auto_in_a_ready(clint_auto_in_a_ready),
    .auto_in_a_valid(clint_auto_in_a_valid),
    .auto_in_a_bits_opcode(clint_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(clint_auto_in_a_bits_size),
    .auto_in_a_bits_source(clint_auto_in_a_bits_source),
    .auto_in_a_bits_address(clint_auto_in_a_bits_address),
    .auto_in_a_bits_mask(clint_auto_in_a_bits_mask),
    .auto_in_a_bits_data(clint_auto_in_a_bits_data),
    .auto_in_d_ready(clint_auto_in_d_ready),
    .auto_in_d_valid(clint_auto_in_d_valid),
    .auto_in_d_bits_opcode(clint_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(clint_auto_in_d_bits_size),
    .auto_in_d_bits_source(clint_auto_in_d_bits_source),
    .auto_in_d_bits_data(clint_auto_in_d_bits_data),
    .io_rtcTick(clint_io_rtcTick),
    .io_covSum(clint_io_covSum)
  );
  IntXbar xbar ( // @[Xbar.scala 30:26]
    .auto_int_in_0(xbar_auto_int_in_0),
    .auto_int_out_0(xbar_auto_int_out_0),
    .io_covSum(xbar_io_covSum)
  );
  IntXbar xbar_1 ( // @[Xbar.scala 30:26]
    .auto_int_in_0(xbar_1_auto_int_in_0),
    .auto_int_out_0(xbar_1_auto_int_out_0),
    .io_covSum(xbar_1_io_covSum)
  );
  IntXbar xbar_2 ( // @[Xbar.scala 30:26]
    .auto_int_in_0(xbar_2_auto_int_in_0),
    .auto_int_out_0(xbar_2_auto_int_out_0),
    .io_covSum(xbar_2_io_covSum)
  );
  BundleBridgeNexus_15 tileHartIdNexusNode ( // @[HasTiles.scala 159:39]
    .auto_out(tileHartIdNexusNode_auto_out),
    .io_covSum(tileHartIdNexusNode_io_covSum)
  );
  IntSyncCrossingSource_4 intsource ( // @[Crossing.scala 26:31]
    .clock(intsource_clock),
    .reset(intsource_reset),
    .auto_in_0(intsource_auto_in_0),
    .auto_in_1(intsource_auto_in_1),
    .auto_out_sync_0(intsource_auto_out_sync_0),
    .auto_out_sync_1(intsource_auto_out_sync_1),
    .io_covSum(intsource_io_covSum)
  );
  IntSyncCrossingSource_1 intsource_1 ( // @[Crossing.scala 26:31]
    .clock(intsource_1_clock),
    .reset(intsource_1_reset),
    .auto_in_0(intsource_1_auto_in_0),
    .auto_out_sync_0(intsource_1_auto_out_sync_0),
    .io_covSum(intsource_1_io_covSum)
  );
  IntSyncCrossingSource_1 intsource_2 ( // @[Crossing.scala 26:31]
    .clock(intsource_2_clock),
    .reset(intsource_2_reset),
    .auto_in_0(intsource_2_auto_in_0),
    .auto_out_sync_0(intsource_2_auto_out_sync_0),
    .io_covSum(intsource_2_io_covSum)
  );
  IntSyncSyncCrossingSink_1 intsink_1 ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_1_auto_in_sync_0),
    .auto_out_0(intsink_1_auto_out_0),
    .io_covSum(intsink_1_io_covSum)
  );
  IntSyncSyncCrossingSink_1 intsink_2 ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_2_auto_in_sync_0),
    .auto_out_0(intsink_2_auto_out_0),
    .io_covSum(intsink_2_io_covSum)
  );
  IntSyncSyncCrossingSink_1 intsink_3 ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_3_auto_in_sync_0),
    .auto_out_0(intsink_3_auto_out_0),
    .io_covSum(intsink_3_io_covSum)
  );
  ClockSinkDomain_1 bootROMDomainWrapper ( // @[BootROM.scala 70:42]
    .auto_bootrom_in_a_ready(bootROMDomainWrapper_auto_bootrom_in_a_ready),
    .auto_bootrom_in_a_valid(bootROMDomainWrapper_auto_bootrom_in_a_valid),
    .auto_bootrom_in_a_bits_size(bootROMDomainWrapper_auto_bootrom_in_a_bits_size),
    .auto_bootrom_in_a_bits_source(bootROMDomainWrapper_auto_bootrom_in_a_bits_source),
    .auto_bootrom_in_a_bits_address(bootROMDomainWrapper_auto_bootrom_in_a_bits_address),
    .auto_bootrom_in_d_ready(bootROMDomainWrapper_auto_bootrom_in_d_ready),
    .auto_bootrom_in_d_valid(bootROMDomainWrapper_auto_bootrom_in_d_valid),
    .auto_bootrom_in_d_bits_size(bootROMDomainWrapper_auto_bootrom_in_d_bits_size),
    .auto_bootrom_in_d_bits_source(bootROMDomainWrapper_auto_bootrom_in_d_bits_source),
    .auto_bootrom_in_d_bits_data(bootROMDomainWrapper_auto_bootrom_in_d_bits_data),
    .io_covSum(bootROMDomainWrapper_io_covSum)
  );
  TLMaskROM maskROM ( // @[MaskROM.scala 66:29]
    .clock(maskROM_clock),
    .reset(maskROM_reset),
    .auto_in_a_ready(maskROM_auto_in_a_ready),
    .auto_in_a_valid(maskROM_auto_in_a_valid),
    .auto_in_a_bits_size(maskROM_auto_in_a_bits_size),
    .auto_in_a_bits_source(maskROM_auto_in_a_bits_source),
    .auto_in_a_bits_address(maskROM_auto_in_a_bits_address),
    .auto_in_d_ready(maskROM_auto_in_d_ready),
    .auto_in_d_valid(maskROM_auto_in_d_valid),
    .auto_in_d_bits_size(maskROM_auto_in_d_bits_size),
    .auto_in_d_bits_source(maskROM_auto_in_d_bits_source),
    .auto_in_d_bits_data(maskROM_auto_in_d_bits_data),
    .io_covSum(maskROM_io_covSum),
    .metaReset(maskROM_metaReset)
  );
  ClockSinkDomain_2 uartClockDomainWrapper ( // @[UART.scala 242:44]
    .auto_uart_0_int_xing_out_sync_0(uartClockDomainWrapper_auto_uart_0_int_xing_out_sync_0),
    .auto_uart_0_control_xing_in_a_ready(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_ready),
    .auto_uart_0_control_xing_in_a_valid(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_valid),
    .auto_uart_0_control_xing_in_a_bits_opcode(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_opcode),
    .auto_uart_0_control_xing_in_a_bits_size(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_size),
    .auto_uart_0_control_xing_in_a_bits_source(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_source),
    .auto_uart_0_control_xing_in_a_bits_address(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_address),
    .auto_uart_0_control_xing_in_a_bits_mask(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_mask),
    .auto_uart_0_control_xing_in_a_bits_data(uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_data),
    .auto_uart_0_control_xing_in_d_ready(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_ready),
    .auto_uart_0_control_xing_in_d_valid(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_valid),
    .auto_uart_0_control_xing_in_d_bits_opcode(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_opcode),
    .auto_uart_0_control_xing_in_d_bits_size(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_size),
    .auto_uart_0_control_xing_in_d_bits_source(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_source),
    .auto_uart_0_control_xing_in_d_bits_data(uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_data),
    .auto_uart_0_io_out_txd(uartClockDomainWrapper_auto_uart_0_io_out_txd),
    .auto_uart_0_io_out_rxd(uartClockDomainWrapper_auto_uart_0_io_out_rxd),
    .auto_clock_in_clock(uartClockDomainWrapper_auto_clock_in_clock),
    .auto_clock_in_reset(uartClockDomainWrapper_auto_clock_in_reset),
    .io_covSum(uartClockDomainWrapper_io_covSum),
    .metaReset(uartClockDomainWrapper_metaReset)
  );
  IntSyncSyncCrossingSink_1 intsink_4 ( // @[Crossing.scala 94:29]
    .auto_in_sync_0(intsink_4_auto_in_sync_0),
    .auto_out_0(intsink_4_auto_out_0),
    .io_covSum(intsink_4_io_covSum)
  );
  MagicDevice magic ( // @[Magic.scala 90:27]
    .clock(magic_clock),
    .reset(magic_reset),
    .auto_in_a_ready(magic_auto_in_a_ready),
    .auto_in_a_valid(magic_auto_in_a_valid),
    .auto_in_a_bits_opcode(magic_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(magic_auto_in_a_bits_size),
    .auto_in_a_bits_source(magic_auto_in_a_bits_source),
    .auto_in_a_bits_address(magic_auto_in_a_bits_address),
    .auto_in_a_bits_mask(magic_auto_in_a_bits_mask),
    .auto_in_d_ready(magic_auto_in_d_ready),
    .auto_in_d_valid(magic_auto_in_d_valid),
    .auto_in_d_bits_opcode(magic_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(magic_auto_in_d_bits_size),
    .auto_in_d_bits_source(magic_auto_in_d_bits_source),
    .auto_in_d_bits_data(magic_auto_in_d_bits_data),
    .io_covSum(magic_io_covSum)
  );
  assign ibus_auto_int_bus_int_out_0 = ibus_int_bus_auto_int_out_0; // @[LazyModule.scala 311:12]
  assign ibus_int_bus_auto_int_in_0 = ibus_auto_int_bus_int_in_0; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_clock =
    subsystem_fbus_subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_reset =
    subsystem_fbus_subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_clockGroup_auto_out_clock = subsystem_fbus_clockGroup_auto_in_member_subsystem_fbus_0_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_clockGroup_auto_out_reset = subsystem_fbus_clockGroup_auto_in_member_subsystem_fbus_0_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_fixedClockNode_auto_out_clock = subsystem_fbus_fixedClockNode_auto_in_clock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_fixedClockNode_auto_out_reset = subsystem_fbus_fixedClockNode_auto_in_reset; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_ready = subsystem_fbus_subsystem_fbus_xbar_auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_d_valid = subsystem_fbus_subsystem_fbus_xbar_auto_out_d_valid; // @[ReadyValidCancel.scala 21:38]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_opcode =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_size =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_source =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_source; // @[Xbar.scala 228:69]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_denied =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_data =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_corrupt =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_valid = subsystem_fbus_subsystem_fbus_xbar_auto_in_a_valid; // @[ReadyValidCancel.scala 21:38]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_opcode =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_param =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_size =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_source =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_source; // @[Xbar.scala 237:55]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_address =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_bufferable =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_modifiable =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_readalloc =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_writealloc =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_privileged =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_secure =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_fetch =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_mask =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_data =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_d_ready = subsystem_fbus_subsystem_fbus_xbar_auto_in_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_ready =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_ready; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_ready =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_ready; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_valid =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_valid; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_bits_id =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_bits_id; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_bits_resp =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_bits_resp; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_ready =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_ready; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_valid =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_valid; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_id =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_id; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_data =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_data; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_resp =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_resp; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_last =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_bits_last; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_auto_bus_xing_out_a_valid = subsystem_fbus_buffer_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_opcode = subsystem_fbus_buffer_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_param = subsystem_fbus_buffer_auto_out_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_size = subsystem_fbus_buffer_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_source = subsystem_fbus_buffer_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_address = subsystem_fbus_buffer_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_bufferable =
    subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_bufferable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_modifiable =
    subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_modifiable; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_readalloc =
    subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_readalloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_writealloc =
    subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_writealloc; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_privileged =
    subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_privileged; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_secure =
    subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_secure; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_fetch =
    subsystem_fbus_buffer_auto_out_a_bits_user_amba_prot_fetch; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_mask = subsystem_fbus_buffer_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_a_bits_data = subsystem_fbus_buffer_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_d_ready = subsystem_fbus_buffer_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_clock =
    subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_reset =
    subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_clockGroup_auto_in_member_subsystem_fbus_0_clock =
    subsystem_fbus_subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_clock; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_clockGroup_auto_in_member_subsystem_fbus_0_reset =
    subsystem_fbus_subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_reset; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_fixedClockNode_auto_in_clock = subsystem_fbus_clockGroup_auto_out_clock; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_fixedClockNode_auto_in_reset = subsystem_fbus_clockGroup_auto_out_reset; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_valid =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_valid; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_opcode =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_param =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_size =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_source =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_address =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_bufferable =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_modifiable =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_readalloc =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_writealloc =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_privileged =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_secure =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_user_amba_prot_fetch =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_mask =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_a_bits_data =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_in_d_ready =
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_ready; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_a_ready = subsystem_fbus_buffer_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_d_valid = subsystem_fbus_buffer_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_opcode = subsystem_fbus_buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_size = subsystem_fbus_buffer_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_source = subsystem_fbus_buffer_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_denied = subsystem_fbus_buffer_auto_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_data = subsystem_fbus_buffer_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_subsystem_fbus_xbar_auto_out_d_bits_corrupt = subsystem_fbus_buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_clock = subsystem_fbus_fixedClockNode_auto_out_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_buffer_reset = subsystem_fbus_fixedClockNode_auto_out_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_buffer_auto_in_a_valid = subsystem_fbus_subsystem_fbus_xbar_auto_out_a_valid; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_opcode = subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_param = subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_param; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_size = subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_source = subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_address = subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_bufferable =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_modifiable =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_readalloc =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_writealloc =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_privileged =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_secure =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_user_amba_prot_fetch =
    subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_mask = subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_a_bits_data = subsystem_fbus_subsystem_fbus_xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_in_d_ready = subsystem_fbus_subsystem_fbus_xbar_auto_out_d_ready; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_buffer_auto_out_a_ready = subsystem_fbus_auto_bus_xing_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_buffer_auto_out_d_valid = subsystem_fbus_auto_bus_xing_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_buffer_auto_out_d_bits_opcode = subsystem_fbus_auto_bus_xing_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_buffer_auto_out_d_bits_size = subsystem_fbus_auto_bus_xing_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_buffer_auto_out_d_bits_source = subsystem_fbus_auto_bus_xing_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_buffer_auto_out_d_bits_denied = subsystem_fbus_auto_bus_xing_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_buffer_auto_out_d_bits_data = subsystem_fbus_auto_bus_xing_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_buffer_auto_out_d_bits_corrupt = subsystem_fbus_auto_bus_xing_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_clock = subsystem_fbus_fixedClockNode_auto_out_clock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_reset = subsystem_fbus_fixedClockNode_auto_out_reset; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_valid =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_valid; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_id =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_id; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_addr =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_addr; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_len =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_len; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_size =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_size; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_burst =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_burst; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_cache =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_cache; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_aw_bits_prot =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_prot; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_valid =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_valid; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_bits_data =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_bits_data; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_bits_strb =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_bits_strb; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_w_bits_last =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_bits_last; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_b_ready =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_ready; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_valid =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_valid; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_id =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_id; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_addr =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_addr; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_len =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_len; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_size =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_size; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_burst =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_burst; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_cache =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_cache; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_ar_bits_prot =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_prot; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_axi4index_in_r_ready =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_ready; // @[LazyModule.scala 309:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_ready =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_a_ready; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_valid =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_d_valid; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_opcode =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_size =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_source =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_denied =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_data =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_bits_corrupt =
    subsystem_fbus_subsystem_fbus_xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign mem_axi4_0_aw_valid = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_aw_bits_id =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_aw_bits_addr =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_aw_bits_len =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_aw_bits_size =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_aw_bits_burst =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_aw_bits_lock =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_lock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_aw_bits_cache =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_aw_bits_prot =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_aw_bits_qos =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_qos; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_w_valid = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_w_bits_data =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_w_bits_strb =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_w_bits_last =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_b_ready = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_valid = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_bits_id =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_bits_addr =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_bits_len =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_bits_size =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_bits_burst =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_bits_lock =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_lock; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_bits_cache =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_cache; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_bits_prot =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_prot; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_ar_bits_qos =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_qos; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign mem_axi4_0_r_ready = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign l2_frontend_bus_axi4_0_aw_ready =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_w_ready =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_b_valid =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_b_bits_id =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_b_bits_resp =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_ar_ready =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_r_valid =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_r_bits_id =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_id; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_r_bits_data =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_r_bits_resp =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_resp; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign l2_frontend_bus_axi4_0_r_bits_last =
    subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_bits_last; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign uart_0_txd = uartClockDomainWrapper_auto_uart_0_io_out_txd; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign ibus_auto_int_bus_int_in_0 = intsink_4_auto_out_0; // @[LazyModule.scala 296:16]
  assign dummyClockGroupSourceNode_clock = clock;
  assign dummyClockGroupSourceNode_reset = reset;
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_valid =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_valid; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_opcode =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_param =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_size =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_source =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_address =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_bufferable =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_modifiable =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_readalloc =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_writealloc =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_privileged =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_secure =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_user_amba_prot_fetch =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_mask =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_bits_data =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_ready =
    tile_prci_domain_auto_tl_master_clock_xing_out_d_ready; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready =
    subsystem_l2_wrapper_auto_coherent_jbar_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid =
    subsystem_fbus_auto_bus_xing_out_a_valid; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode =
    subsystem_fbus_auto_bus_xing_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param =
    subsystem_fbus_auto_bus_xing_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size =
    subsystem_fbus_auto_bus_xing_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source =
    subsystem_fbus_auto_bus_xing_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address =
    subsystem_fbus_auto_bus_xing_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_bufferable =
    subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_modifiable =
    subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_readalloc =
    subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_writealloc =
    subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_privileged =
    subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_secure =
    subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_user_amba_prot_fetch =
    subsystem_fbus_auto_bus_xing_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask =
    subsystem_fbus_auto_bus_xing_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data =
    subsystem_fbus_auto_bus_xing_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready =
    subsystem_fbus_auto_bus_xing_out_d_ready; // @[LazyModule.scala 296:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready =
    subsystem_cbus_auto_bus_xing_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid =
    subsystem_cbus_auto_bus_xing_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode =
    subsystem_cbus_auto_bus_xing_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size =
    subsystem_cbus_auto_bus_xing_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source =
    subsystem_cbus_auto_bus_xing_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied =
    subsystem_cbus_auto_bus_xing_in_d_bits_denied; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data =
    subsystem_cbus_auto_bus_xing_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt =
    subsystem_cbus_auto_bus_xing_in_d_bits_corrupt; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_clock; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_reset; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_clock; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_reset; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_clock; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_reset; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_clock; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_reset; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_clock; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_reset; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_clock; // @[LazyModule.scala 298:16]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_reset; // @[LazyModule.scala 298:16]
  assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_ready =
    uartClockDomainWrapper_auto_uart_0_control_xing_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_valid =
    uartClockDomainWrapper_auto_uart_0_control_xing_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_opcode =
    uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_size =
    uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_source =
    uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_bits_data =
    uartClockDomainWrapper_auto_uart_0_control_xing_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock =
    subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset =
    subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_bus_xing_in_a_valid =
    subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_valid; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_bus_xing_in_a_bits_opcode =
    subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_bus_xing_in_a_bits_param =
    subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_bus_xing_in_a_bits_size =
    subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_bus_xing_in_a_bits_source =
    subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_bus_xing_in_a_bits_address =
    subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_bus_xing_in_a_bits_mask =
    subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_bus_xing_in_a_bits_data =
    subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_pbus_auto_bus_xing_in_d_ready =
    subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_ready; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_valid =
    l2_frontend_bus_axi4_0_aw_valid; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_id =
    l2_frontend_bus_axi4_0_aw_bits_id; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_addr =
    l2_frontend_bus_axi4_0_aw_bits_addr; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_len =
    l2_frontend_bus_axi4_0_aw_bits_len; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_size =
    l2_frontend_bus_axi4_0_aw_bits_size; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_burst =
    l2_frontend_bus_axi4_0_aw_bits_burst; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_cache =
    l2_frontend_bus_axi4_0_aw_bits_cache; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_aw_bits_prot =
    l2_frontend_bus_axi4_0_aw_bits_prot; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_valid =
    l2_frontend_bus_axi4_0_w_valid; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_bits_data =
    l2_frontend_bus_axi4_0_w_bits_data; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_bits_strb =
    l2_frontend_bus_axi4_0_w_bits_strb; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_w_bits_last =
    l2_frontend_bus_axi4_0_w_bits_last; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_b_ready =
    l2_frontend_bus_axi4_0_b_ready; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_valid =
    l2_frontend_bus_axi4_0_ar_valid; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_id =
    l2_frontend_bus_axi4_0_ar_bits_id; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_addr =
    l2_frontend_bus_axi4_0_ar_bits_addr; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_len =
    l2_frontend_bus_axi4_0_ar_bits_len; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_size =
    l2_frontend_bus_axi4_0_ar_bits_size; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_burst =
    l2_frontend_bus_axi4_0_ar_bits_burst; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_cache =
    l2_frontend_bus_axi4_0_ar_bits_cache; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_ar_bits_prot =
    l2_frontend_bus_axi4_0_ar_bits_prot; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_coupler_from_port_named_slave_port_axi4_axi4index_in_r_ready =
    l2_frontend_bus_axi4_0_r_ready; // @[Nodes.scala 1207:84 1630:60]
  assign subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset; // @[LazyModule.scala 298:16]
  assign subsystem_fbus_auto_bus_xing_out_a_ready =
    subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_d_valid =
    subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_d_bits_opcode =
    subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_d_bits_size =
    subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_d_bits_source =
    subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_d_bits_denied =
    subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_d_bits_data =
    subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_fbus_auto_bus_xing_out_d_bits_corrupt =
    subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_ready = magic_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_valid = magic_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_opcode = magic_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_size = magic_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_source = magic_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_bits_data = magic_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_ready = maskROM_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_valid = maskROM_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_bits_size = maskROM_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_bits_source = maskROM_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_bits_data = maskROM_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_ready = bootROMDomainWrapper_auto_bootrom_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_valid = bootROMDomainWrapper_auto_bootrom_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_size =
    bootROMDomainWrapper_auto_bootrom_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_source =
    bootROMDomainWrapper_auto_bootrom_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_data =
    bootROMDomainWrapper_auto_bootrom_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_ready = clint_auto_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_valid = clint_auto_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_opcode = clint_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_size = clint_auto_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_source = clint_auto_in_d_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_bits_data = clint_auto_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_ready = plicDomainWrapper_auto_plic_in_a_ready; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_valid = plicDomainWrapper_auto_plic_in_d_valid; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_opcode = plicDomainWrapper_auto_plic_in_d_bits_opcode
    ; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_size = plicDomainWrapper_auto_plic_in_d_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_source = plicDomainWrapper_auto_plic_in_d_bits_source
    ; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_bits_data = plicDomainWrapper_auto_plic_in_d_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_a_ready =
    subsystem_pbus_auto_bus_xing_in_a_ready; // @[LazyModule.scala 296:16]
  assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_valid =
    subsystem_pbus_auto_bus_xing_in_d_valid; // @[LazyModule.scala 296:16]
  assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_opcode =
    subsystem_pbus_auto_bus_xing_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_size =
    subsystem_pbus_auto_bus_xing_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_source =
    subsystem_pbus_auto_bus_xing_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_denied =
    subsystem_pbus_auto_bus_xing_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_data =
    subsystem_pbus_auto_bus_xing_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_cbus_auto_coupler_to_bus_named_subsystem_pbus_bus_xing_out_d_bits_corrupt =
    subsystem_pbus_auto_bus_xing_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_bus_xing_in_a_valid =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_opcode =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_param =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_size =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_source =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_address =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_mask =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_data =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_cbus_auto_bus_xing_in_d_ready =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready; // @[LazyModule.scala 298:16]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready = mem_axi4_0_aw_ready; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready = mem_axi4_0_w_ready; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid = mem_axi4_0_b_valid; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id = mem_axi4_0_b_bits_id; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp =
    mem_axi4_0_b_bits_resp; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready = mem_axi4_0_ar_ready; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid = mem_axi4_0_r_valid; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id = mem_axi4_0_r_bits_id; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data =
    mem_axi4_0_r_bits_data; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp =
    mem_axi4_0_r_bits_resp; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last =
    mem_axi4_0_r_bits_last; // @[Nodes.scala 1210:84 1694:56]
  assign subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock =
    subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset =
    subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_valid =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_opcode =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_size =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_source =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_address =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_bufferable =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_modifiable =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_readalloc =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_writealloc =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_privileged =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_secure =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_user_amba_prot_fetch =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_mask =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_data =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_mbus_auto_bus_xing_in_d_ready =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready; // @[LazyModule.scala 296:16]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready =
    subsystem_mbus_auto_bus_xing_in_a_ready; // @[LazyModule.scala 296:16]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid =
    subsystem_mbus_auto_bus_xing_in_d_valid; // @[LazyModule.scala 296:16]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode =
    subsystem_mbus_auto_bus_xing_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size =
    subsystem_mbus_auto_bus_xing_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source =
    subsystem_mbus_auto_bus_xing_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied =
    subsystem_mbus_auto_bus_xing_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data =
    subsystem_mbus_auto_bus_xing_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt =
    subsystem_mbus_auto_bus_xing_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_valid =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_opcode =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_size =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_source =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_address =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_bufferable =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_bufferable; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_modifiable =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_modifiable; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_readalloc =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_readalloc; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_writealloc =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_writealloc; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_privileged =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_privileged; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_secure =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_secure; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_user_amba_prot_fetch =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_user_amba_prot_fetch; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_mask =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_data =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_d_ready =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock; // @[LazyModule.scala 298:16]
  assign subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset; // @[LazyModule.scala 298:16]
  assign tile_prci_domain_auto_tile_reset_domain_cva6_tile_hartid_in = tileHartIdNexusNode_auto_out; // @[LazyModule.scala 296:16]
  assign tile_prci_domain_auto_int_in_clock_xing_in_2_sync_0 = intsource_2_auto_out_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tile_prci_domain_auto_int_in_clock_xing_in_1_sync_0 = intsource_1_auto_out_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tile_prci_domain_auto_int_in_clock_xing_in_0_sync_0 = intsource_auto_out_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tile_prci_domain_auto_int_in_clock_xing_in_0_sync_1 = intsource_auto_out_sync_1; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_a_ready =
    subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_a_ready; // @[LazyModule.scala 296:16]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_valid =
    subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_valid; // @[LazyModule.scala 296:16]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_opcode =
    subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_size =
    subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_size; // @[LazyModule.scala 296:16]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_source =
    subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_source; // @[LazyModule.scala 296:16]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_denied =
    subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_denied; // @[LazyModule.scala 296:16]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_data =
    subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_data; // @[LazyModule.scala 296:16]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_corrupt =
    subsystem_sbus_auto_coupler_from_cva6_tile_tl_master_clock_xing_in_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign tile_prci_domain_auto_tap_clock_in_clock = subsystem_sbus_auto_fixedClockNode_out_1_clock; // @[LazyModule.scala 298:16]
  assign tile_prci_domain_auto_tap_clock_in_reset = subsystem_sbus_auto_fixedClockNode_out_1_reset; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_plic_int_in_0 = ibus_auto_int_bus_int_out_0; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_plic_in_a_valid = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_valid; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_plic_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_opcode
    ; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_plic_in_a_bits_size = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_plic_in_a_bits_source = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_source
    ; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_plic_in_a_bits_address =
    subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_plic_in_a_bits_mask = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_plic_in_a_bits_data = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_plic_in_d_ready = subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_ready; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_clock_in_clock = subsystem_cbus_auto_fixedClockNode_out_0_clock; // @[LazyModule.scala 298:16]
  assign plicDomainWrapper_auto_clock_in_reset = subsystem_cbus_auto_fixedClockNode_out_0_reset; // @[LazyModule.scala 298:16]
  assign clint_clock = subsystem_cbus_clock; // @[CLINT.scala 115:26]
  assign clint_reset = subsystem_cbus_reset; // @[CLINT.scala 116:26]
  assign clint_auto_in_a_valid = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_valid; // @[LazyModule.scala 298:16]
  assign clint_auto_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign clint_auto_in_a_bits_size = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign clint_auto_in_a_bits_source = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign clint_auto_in_a_bits_address = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign clint_auto_in_a_bits_mask = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign clint_auto_in_a_bits_data = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign clint_auto_in_d_ready = subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_ready; // @[LazyModule.scala 298:16]
  assign clint_io_rtcTick = int_rtc_tick_value == 7'h63; // @[Counter.scala 74:24]
  assign xbar_auto_int_in_0 = intsink_1_auto_out_0; // @[LazyModule.scala 296:16]
  assign xbar_1_auto_int_in_0 = intsink_2_auto_out_0; // @[LazyModule.scala 296:16]
  assign xbar_2_auto_int_in_0 = intsink_3_auto_out_0; // @[LazyModule.scala 296:16]
  assign intsource_clock = clock;
  assign intsource_reset = reset;
  assign intsource_auto_in_0 = clint_auto_int_out_0; // @[LazyModule.scala 298:16]
  assign intsource_auto_in_1 = clint_auto_int_out_1; // @[LazyModule.scala 298:16]
  assign intsource_1_clock = clock;
  assign intsource_1_reset = reset;
  assign intsource_1_auto_in_0 = plicDomainWrapper_auto_plic_int_out_0_0; // @[LazyModule.scala 298:16]
  assign intsource_2_clock = clock;
  assign intsource_2_reset = reset;
  assign intsource_2_auto_in_0 = plicDomainWrapper_auto_plic_int_out_1_0; // @[LazyModule.scala 298:16]
  assign intsink_1_auto_in_sync_0 = tile_prci_domain_auto_int_out_clock_xing_out_0_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign intsink_2_auto_in_sync_0 = tile_prci_domain_auto_int_out_clock_xing_out_1_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign intsink_3_auto_in_sync_0 = tile_prci_domain_auto_int_out_clock_xing_out_2_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign bootROMDomainWrapper_auto_bootrom_in_a_valid = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid; // @[LazyModule.scala 298:16]
  assign bootROMDomainWrapper_auto_bootrom_in_a_bits_size =
    subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign bootROMDomainWrapper_auto_bootrom_in_a_bits_source =
    subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign bootROMDomainWrapper_auto_bootrom_in_a_bits_address =
    subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign bootROMDomainWrapper_auto_bootrom_in_d_ready = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready; // @[LazyModule.scala 298:16]
  assign maskROM_clock = subsystem_cbus_clock; // @[MaskROM.scala 70:41]
  assign maskROM_reset = subsystem_cbus_reset; // @[MaskROM.scala 71:41]
  assign maskROM_auto_in_a_valid = subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_valid; // @[LazyModule.scala 298:16]
  assign maskROM_auto_in_a_bits_size = subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign maskROM_auto_in_a_bits_source = subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign maskROM_auto_in_a_bits_address = subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign maskROM_auto_in_d_ready = subsystem_cbus_auto_coupler_to_MaskROM_fragmenter_out_d_ready; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_valid =
    subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_valid; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_opcode =
    subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_size =
    subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_source =
    subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_address =
    subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_mask =
    subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_uart_0_control_xing_in_a_bits_data =
    subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_a_bits_data; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_uart_0_control_xing_in_d_ready =
    subsystem_pbus_auto_coupler_to_device_named_uart_0_control_xing_out_d_ready; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_uart_0_io_out_rxd = uart_0_rxd; // @[Nodes.scala 1210:84 BundleBridge.scala 54:8]
  assign uartClockDomainWrapper_auto_clock_in_clock = subsystem_pbus_auto_fixedClockNode_out_clock; // @[LazyModule.scala 298:16]
  assign uartClockDomainWrapper_auto_clock_in_reset = subsystem_pbus_auto_fixedClockNode_out_reset; // @[LazyModule.scala 298:16]
  assign intsink_4_auto_in_sync_0 = uartClockDomainWrapper_auto_uart_0_int_xing_out_sync_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign magic_clock = clock;
  assign magic_reset = reset;
  assign magic_auto_in_a_valid = subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_valid; // @[LazyModule.scala 298:16]
  assign magic_auto_in_a_bits_opcode = subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_opcode; // @[LazyModule.scala 298:16]
  assign magic_auto_in_a_bits_size = subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_size; // @[LazyModule.scala 298:16]
  assign magic_auto_in_a_bits_source = subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_source; // @[LazyModule.scala 298:16]
  assign magic_auto_in_a_bits_address = subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_address; // @[LazyModule.scala 298:16]
  assign magic_auto_in_a_bits_mask = subsystem_cbus_auto_coupler_to_magic_fragmenter_out_a_bits_mask; // @[LazyModule.scala 298:16]
  assign magic_auto_in_d_ready = subsystem_cbus_auto_coupler_to_magic_fragmenter_out_d_ready; // @[LazyModule.scala 298:16]
  assign StarshipASICTop_covSum = 30'h0;
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_sum = StarshipASICTop_covSum +
    subsystem_fbus_coupler_from_port_named_slave_port_axi4_io_covSum;
  assign ibus_int_bus_sum = subsystem_fbus_coupler_from_port_named_slave_port_axi4_sum + ibus_int_bus_io_covSum;
  assign intsink_2_sum = ibus_int_bus_sum + intsink_2_io_covSum;
  assign subsystem_fbus_buffer_sum = intsink_2_sum + subsystem_fbus_buffer_io_covSum;
  assign subsystem_l2_wrapper_sum = subsystem_fbus_buffer_sum + subsystem_l2_wrapper_io_covSum;
  assign tile_prci_domain_sum = subsystem_l2_wrapper_sum + tile_prci_domain_io_covSum;
  assign maskROM_sum = tile_prci_domain_sum + maskROM_io_covSum;
  assign subsystem_sbus_sum = maskROM_sum + subsystem_sbus_io_covSum;
  assign subsystem_cbus_sum = subsystem_sbus_sum + subsystem_cbus_io_covSum;
  assign bootROMDomainWrapper_sum = subsystem_cbus_sum + bootROMDomainWrapper_io_covSum;
  assign xbar_1_sum = bootROMDomainWrapper_sum + xbar_1_io_covSum;
  assign intsink_1_sum = xbar_1_sum + intsink_1_io_covSum;
  assign uartClockDomainWrapper_sum = intsink_1_sum + uartClockDomainWrapper_io_covSum;
  assign intsource_1_sum = uartClockDomainWrapper_sum + intsource_1_io_covSum;
  assign tileHartIdNexusNode_sum = intsource_1_sum + tileHartIdNexusNode_io_covSum;
  assign dummyClockGroupSourceNode_sum = tileHartIdNexusNode_sum + dummyClockGroupSourceNode_io_covSum;
  assign magic_sum = dummyClockGroupSourceNode_sum + magic_io_covSum;
  assign subsystem_pbus_sum = magic_sum + subsystem_pbus_io_covSum;
  assign xbar_sum = subsystem_pbus_sum + xbar_io_covSum;
  assign xbar_2_sum = xbar_sum + xbar_2_io_covSum;
  assign subsystem_mbus_sum = xbar_2_sum + subsystem_mbus_io_covSum;
  assign plicDomainWrapper_sum = subsystem_mbus_sum + plicDomainWrapper_io_covSum;
  assign intsource_sum = plicDomainWrapper_sum + intsource_io_covSum;
  assign intsink_4_sum = intsource_sum + intsink_4_io_covSum;
  assign clint_sum = intsink_4_sum + clint_io_covSum;
  assign intsource_2_sum = clint_sum + intsource_2_io_covSum;
  assign intsink_3_sum = intsource_2_sum + intsink_3_io_covSum;
  assign io_covSum = intsink_3_sum;
  assign subsystem_fbus_coupler_from_port_named_slave_port_axi4_metaReset = metaReset;
  assign subsystem_l2_wrapper_metaReset = metaReset;
  assign tile_prci_domain_metaReset = metaReset;
  assign maskROM_metaReset = metaReset;
  assign subsystem_sbus_metaReset = metaReset;
  assign subsystem_cbus_metaReset = metaReset;
  assign uartClockDomainWrapper_metaReset = metaReset;
  assign subsystem_pbus_metaReset = metaReset;
  assign subsystem_mbus_metaReset = metaReset;
  assign plicDomainWrapper_metaReset = metaReset;
  always @(posedge subsystem_pbus_clock) begin
    if (subsystem_pbus_reset) begin // @[Counter.scala 62:40]
      int_rtc_tick_value <= 7'h0; // @[Counter.scala 62:40]
    end else if (int_rtc_tick_wrap_wrap) begin
      int_rtc_tick_value <= 7'h0;
    end else begin
      int_rtc_tick_value <= _int_rtc_tick_wrap_value_T_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  int_rtc_tick_value = _RAND_0[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
